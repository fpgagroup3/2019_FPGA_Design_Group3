module	dense1(
	input clk,
	input rst_n,
	input [256*16-1:0] d1_input,
	output reg [4*16-1:0] d1_output
);


reg [15:0] d1_input_r [0:255];

reg [31:0] temp_mult [0:1023];
reg [15:0] temp_add [0:3];
reg [4:0] counter;
reg [15:0] a,b [0:63];
wire [15:0] bias [0:3];

wire [31:0] mult [0:63];

integer i, j;

assign bias[0] = 16'd346;
assign bias[1] = 16'd344; 
assign bias[2] = 16'd33106; 
assign bias[3] = 16'd33106;

assign mult[0]  = a[0] * b[0];
assign mult[1]  = a[1] * b[1];
assign mult[2]  = a[2] * b[2];
assign mult[3]  = a[3] * b[3];
assign mult[4]  = a[4] * b[4];
assign mult[5]  = a[5] * b[5];
assign mult[6]  = a[6] * b[6];
assign mult[7]  = a[7] * b[7];
assign mult[8]  = a[8] * b[8];
assign mult[9]  = a[9] * b[9];
assign mult[10] = a[10] * b[10];
assign mult[11] = a[11] * b[11];
assign mult[12] = a[12] * b[12];
assign mult[13] = a[13] * b[13];
assign mult[14] = a[14] * b[14];
assign mult[15] = a[15] * b[15];
assign mult[16] = a[16] * b[16];
assign mult[17] = a[17] * b[17];
assign mult[18] = a[18] * b[18];
assign mult[19] = a[19] * b[19];
assign mult[20] = a[20] * b[20];
assign mult[21] = a[21] * b[21];
assign mult[22] = a[22] * b[22];
assign mult[23] = a[23] * b[23];
assign mult[24] = a[24] * b[24];
assign mult[25] = a[25] * b[25];
assign mult[26] = a[26] * b[26];
assign mult[27] = a[27] * b[27];
assign mult[28] = a[28] * b[28];
assign mult[29] = a[29] * b[29];
assign mult[30] = a[30] * b[30];
assign mult[31] = a[31] * b[31];
assign mult[32] = a[32] * b[32];
assign mult[33] = a[33] * b[33];
assign mult[34] = a[34] * b[34];
assign mult[35] = a[35] * b[35];
assign mult[36] = a[36] * b[36];
assign mult[37] = a[37] * b[37];
assign mult[38] = a[38] * b[38];
assign mult[39] = a[39] * b[39];
assign mult[40] = a[40] * b[40];
assign mult[41] = a[41] * b[41];
assign mult[42] = a[42] * b[42];
assign mult[43] = a[43] * b[43];
assign mult[44] = a[44] * b[44];
assign mult[45] = a[45] * b[45];
assign mult[46] = a[46] * b[46];
assign mult[47] = a[47] * b[47];
assign mult[48] = a[48] * b[48];
assign mult[49] = a[49] * b[49];
assign mult[50] = a[50] * b[50];
assign mult[51] = a[51] * b[51];
assign mult[52] = a[52] * b[52];
assign mult[53] = a[53] * b[53];
assign mult[54] = a[54] * b[54];
assign mult[55] = a[55] * b[55];
assign mult[56] = a[56] * b[56];
assign mult[57] = a[57] * b[57];
assign mult[58] = a[58] * b[58];
assign mult[59] = a[59] * b[59];
assign mult[60] = a[60] * b[60];
assign mult[61] = a[61] * b[61];
assign mult[62] = a[62] * b[62];
assign mult[63] = a[63] * b[63];


always @(*) begin
	if(!rst_n) begin
		for(j = 0; j < 256; j = j+1) begin
			d1_input_r[j] = 16'd0;
		end
	end
	else begin
		for(j = 0; j < 256; j = j+1) begin
			d1_input_r[j] = d1_input[((16*(j+1))-1) -: 16];
		end
	end
end

always @(*) begin
	case(counter)
		5'd1: begin
			b[0]  =  d1_input_r[0];
			b[1]  =  d1_input_r[1];
			b[2]  =  d1_input_r[2];
			b[3]  =  d1_input_r[3];
			b[4]  =  d1_input_r[4];
			b[5]  =  d1_input_r[5];
			b[6]  =  d1_input_r[6];
			b[7]  =  d1_input_r[7];
			b[8]  =  d1_input_r[8];
			b[9]  =  d1_input_r[9];
			b[10] =  d1_input_r[10];
			b[11] =  d1_input_r[11];
			b[12] =  d1_input_r[12];
			b[13] =  d1_input_r[13];
			b[14] =  d1_input_r[14];
			b[15] =  d1_input_r[15];
			b[16] =  d1_input_r[16];
			b[17] =  d1_input_r[17];
			b[18] =  d1_input_r[18];
			b[19] =  d1_input_r[19];
			b[20] =  d1_input_r[20];
			b[21] =  d1_input_r[21];
			b[22] =  d1_input_r[22];
			b[23] =  d1_input_r[23];
			b[24] =  d1_input_r[24];
			b[25] =  d1_input_r[25];
			b[26] =  d1_input_r[26];
			b[27] =  d1_input_r[27];
			b[28] =  d1_input_r[28];
			b[29] =  d1_input_r[29];
			b[30] =  d1_input_r[30];
			b[31] =  d1_input_r[31];
			b[32] =  d1_input_r[32];
			b[33] =  d1_input_r[33];
			b[34] =  d1_input_r[34];
			b[35] =  d1_input_r[35];
			b[36] =  d1_input_r[36];
			b[37] =  d1_input_r[37];
			b[38] =  d1_input_r[38];
			b[39] =  d1_input_r[39];
			b[40] =  d1_input_r[40];
			b[41] =  d1_input_r[41];
			b[42] =  d1_input_r[42];
			b[43] =  d1_input_r[43];
			b[44] =  d1_input_r[44];
			b[45] =  d1_input_r[45];
			b[46] =  d1_input_r[46];
			b[47] =  d1_input_r[47];
			b[48] =  d1_input_r[48];
			b[49] =  d1_input_r[49];
			b[50] =  d1_input_r[50];
			b[51] =  d1_input_r[51];
			b[52] =  d1_input_r[52];
			b[53] =  d1_input_r[53];
			b[54] =  d1_input_r[54];
			b[55] =  d1_input_r[55];
			b[56] =  d1_input_r[56];
			b[57] =  d1_input_r[57];
			b[58] =  d1_input_r[58];
			b[59] =  d1_input_r[59];
			b[60] =  d1_input_r[60];
			b[61] =  d1_input_r[61];
			b[62] =  d1_input_r[62];
			b[63] =  d1_input_r[63];
			a[0]  =  16'd33087;
			a[1]  =  16'd198  ;
			a[2]  =  16'd34748;
			a[3]  =  16'd2210 ;
			a[4]  =  16'd1852 ;
			a[5]  =  16'd1435 ;
			a[6]  =  16'd157  ;
			a[7]  =  16'd1119 ;
			a[8]  =  16'd1120 ;
			a[9]  =  16'd986  ;
			a[10] =  16'd1497 ;
			a[11] =  16'd993  ;
			a[12] =  16'd35132;
			a[13] =  16'd2385 ;
			a[14] =  16'd2952 ;
			a[15] =  16'd35274;
			a[16] =  16'd33781;
			a[17] =  16'd1008 ;
			a[18] =  16'd560  ;
			a[19] =  16'd1522 ;
			a[20] =  16'd33187;
			a[21] =  16'd490  ;
			a[22] =  16'd581  ;
			a[23] =  16'd33711;
			a[24] =  16'd32952;
			a[25] =  16'd1612 ;
			a[26] =  16'd948  ;
			a[27] =  16'd94   ;
			a[28] =  16'd32906;
			a[29] =  16'd34931;
			a[30] =  16'd33268;
			a[31] =  16'd33834;
			a[32] =  16'd138  ;
			a[33] =  16'd33917;
			a[34] =  16'd1104 ;
			a[35] =  16'd34255;
			a[36] =  16'd34349;
			a[37] =  16'd33242;
			a[38] =  16'd33852;
			a[39] =  16'd717  ;
			a[40] =  16'd1312 ;
			a[41] =  16'd35246;
			a[42] =  16'd2851 ;
			a[43] =  16'd36   ;
			a[44] =  16'd35195;
			a[45] =  16'd35256;
			a[46] =  16'd35134;
			a[47] =  16'd1111 ;
			a[48] =  16'd816  ;
			a[49] =  16'd1649 ;
			a[50] =  16'd33560;
			a[51] =  16'd33982;
			a[52] =  16'd1348 ;
			a[53] =  16'd1352 ;
			a[54] =  16'd870  ;
			a[55] =  16'd1299 ;
			a[56] =  16'd1142 ;
			a[57] =  16'd33779;
			a[58] =  16'd34197;
			a[59] =  16'd174  ;
			a[60] =  16'd2467 ;
			a[61] =  16'd787  ;
			a[62] =  16'd309  ;
			a[63] =  16'd33043;
			temp_mult[0]  = mult[0] ;
			temp_mult[1]  = mult[1] ;
			temp_mult[2]  = mult[2] ;
			temp_mult[3]  = mult[3] ;
			temp_mult[4]  = mult[4] ;
			temp_mult[5]  = mult[5] ;
			temp_mult[6]  = mult[6] ;
			temp_mult[7]  = mult[7] ;
			temp_mult[8]  = mult[8] ;
			temp_mult[9]  = mult[9] ;
			temp_mult[10] = mult[10];
			temp_mult[11] = mult[11];
			temp_mult[12] = mult[12];
			temp_mult[13] = mult[13];
			temp_mult[14] = mult[14];
			temp_mult[15] = mult[15];
			temp_mult[16] = mult[16];
			temp_mult[17] = mult[17];
			temp_mult[18] = mult[18];
			temp_mult[19] = mult[19];
			temp_mult[20] = mult[20];
			temp_mult[21] = mult[21];
			temp_mult[22] = mult[22];
			temp_mult[23] = mult[23];
			temp_mult[24] = mult[24];
			temp_mult[25] = mult[25];
			temp_mult[26] = mult[26];
			temp_mult[27] = mult[27];
			temp_mult[28] = mult[28];
			temp_mult[29] = mult[29];
			temp_mult[30] = mult[30];
			temp_mult[31] = mult[31];
			temp_mult[32] = mult[32];
			temp_mult[33] = mult[33];
			temp_mult[34] = mult[34];
			temp_mult[35] = mult[35];
			temp_mult[36] = mult[36];
			temp_mult[37] = mult[37];
			temp_mult[38] = mult[38];
			temp_mult[39] = mult[39];
			temp_mult[40] = mult[40];
			temp_mult[41] = mult[41];
			temp_mult[42] = mult[42];
			temp_mult[43] = mult[43];
			temp_mult[44] = mult[44];
			temp_mult[45] = mult[45];
			temp_mult[46] = mult[46];
			temp_mult[47] = mult[47];
			temp_mult[48] = mult[48];
			temp_mult[49] = mult[49];
			temp_mult[50] = mult[50];
			temp_mult[51] = mult[51];
			temp_mult[52] = mult[52];
			temp_mult[53] = mult[53];
			temp_mult[54] = mult[54];
			temp_mult[55] = mult[55];
			temp_mult[56] = mult[56];
			temp_mult[57] = mult[57];
			temp_mult[58] = mult[58];
			temp_mult[59] = mult[59];
			temp_mult[60] = mult[60];
			temp_mult[61] = mult[61];
			temp_mult[62] = mult[62];
			temp_mult[63] = mult[63];
		end
		5'd2: begin
			b[0]  = d1_input_r[64];
			b[1]  = d1_input_r[65];
			b[2]  = d1_input_r[66];
			b[3]  = d1_input_r[67];
			b[4]  = d1_input_r[68];
			b[5]  = d1_input_r[69];
			b[6]  = d1_input_r[70];
			b[7]  = d1_input_r[71];
			b[8]  = d1_input_r[72];
			b[9]  = d1_input_r[73];
			b[10] = d1_input_r[74];
			b[11] = d1_input_r[75];
			b[12] = d1_input_r[76];
			b[13] = d1_input_r[77];
			b[14] = d1_input_r[78];
			b[15] = d1_input_r[79];
			b[16] = d1_input_r[80];
			b[17] = d1_input_r[81];
			b[18] = d1_input_r[82];
			b[19] = d1_input_r[83];
			b[20] = d1_input_r[84];
			b[21] = d1_input_r[85];
			b[22] = d1_input_r[86];
			b[23] = d1_input_r[87];
			b[24] = d1_input_r[88];
			b[25] = d1_input_r[89];
			b[26] = d1_input_r[90];
			b[27] = d1_input_r[91];
			b[28] = d1_input_r[92];
			b[29] = d1_input_r[93];
			b[30] = d1_input_r[94];
			b[31] = d1_input_r[95];
			b[32] = d1_input_r[96];
			b[33] = d1_input_r[97];
			b[34] = d1_input_r[98];
			b[35] = d1_input_r[99];
			b[36] = d1_input_r[100];
			b[37] = d1_input_r[101];
			b[38] = d1_input_r[102];
			b[39] = d1_input_r[103];
			b[40] = d1_input_r[104];
			b[41] = d1_input_r[105];
			b[42] = d1_input_r[106];
			b[43] = d1_input_r[107];
			b[44] = d1_input_r[108];
			b[45] = d1_input_r[109];
			b[46] = d1_input_r[110];
			b[47] = d1_input_r[111];
			b[48] = d1_input_r[112];
			b[49] = d1_input_r[113];
			b[50] = d1_input_r[114];
			b[51] = d1_input_r[115];
			b[52] = d1_input_r[116];
			b[53] = d1_input_r[117];
			b[54] = d1_input_r[118];
			b[55] = d1_input_r[119];
			b[56] = d1_input_r[120];
			b[57] = d1_input_r[121];
			b[58] = d1_input_r[122];
			b[59] = d1_input_r[123];
			b[60] = d1_input_r[124];
			b[61] = d1_input_r[125];
			b[62] = d1_input_r[126];
			b[63] = d1_input_r[127];
			a[0]  = 16'd33899;
			a[1]  = 16'd32983;
			a[2]  = 16'd2133 ;
			a[3]  = 16'd1803 ;
			a[4]  = 16'd1557 ;
			a[5]  = 16'd169  ;
			a[6]  = 16'd1054 ;
			a[7]  = 16'd1449 ;
			a[8]  = 16'd32910;
			a[9]  = 16'd34527;
			a[10] = 16'd1212 ;
			a[11] = 16'd1618 ;
			a[12] = 16'd1457 ;
			a[13] = 16'd563  ;
			a[14] = 16'd33332;
			a[15] = 16'd32956;
			a[16] = 16'd1281 ;
			a[17] = 16'd33648;
			a[18] = 16'd1407 ;
			a[19] = 16'd34453;
			a[20] = 16'd35037;
			a[21] = 16'd900  ;
			a[22] = 16'd120  ;
			a[23] = 16'd35796;
			a[24] = 16'd34609;
			a[25] = 16'd35377;
			a[26] = 16'd1416 ;
			a[27] = 16'd34359;
			a[28] = 16'd2394 ;
			a[29] = 16'd698  ;
			a[30] = 16'd32824;
			a[31] = 16'd33476;
			a[32] = 16'd2785 ;
			a[33] = 16'd33356;
			a[34] = 16'd2651 ;
			a[35] = 16'd33599;
			a[36] = 16'd33773;
			a[37] = 16'd726  ;
			a[38] = 16'd1019 ;
			a[39] = 16'd83   ;
			a[40] = 16'd34379;
			a[41] = 16'd34386;
			a[42] = 16'd34448;
			a[43] = 16'd33480;
			a[44] = 16'd881  ;
			a[45] = 16'd34240;
			a[46] = 16'd1850 ;
			a[47] = 16'd33793;
			a[48] = 16'd33106;
			a[49] = 16'd2276 ;
			a[50] = 16'd33897;
			a[51] = 16'd411  ;
			a[52] = 16'd1711 ;
			a[53] = 16'd2660 ;
			a[54] = 16'd33161;
			a[55] = 16'd2370 ;
			a[56] = 16'd458  ;
			a[57] = 16'd33115;
			a[58] = 16'd34893;
			a[59] = 16'd33368;
			a[60] = 16'd2285 ;
			a[61] = 16'd415  ;
			a[62] = 16'd656  ;
			a[63] = 16'd147  ;
			temp_mult[64] = mult[0] ;
			temp_mult[65] = mult[1] ;
			temp_mult[66] = mult[2] ;
			temp_mult[67] = mult[3] ;
			temp_mult[68] = mult[4] ;
			temp_mult[69] = mult[5] ;
			temp_mult[70] = mult[6] ;
			temp_mult[71] = mult[7] ;
			temp_mult[72] = mult[8] ;
			temp_mult[73] = mult[9] ;
			temp_mult[74] = mult[10];
			temp_mult[75] = mult[11];
			temp_mult[76] = mult[12];
			temp_mult[77] = mult[13];
			temp_mult[78] = mult[14];
			temp_mult[79] = mult[15];
			temp_mult[80] = mult[16];
			temp_mult[81] = mult[17];
			temp_mult[82] = mult[18];
			temp_mult[83] = mult[19];
			temp_mult[84] = mult[20];
			temp_mult[85] = mult[21];
			temp_mult[86] = mult[22];
			temp_mult[87] = mult[23];
			temp_mult[88] = mult[24];
			temp_mult[89] = mult[25];
			temp_mult[90] = mult[26];
			temp_mult[91] = mult[27];
			temp_mult[92] = mult[28];
			temp_mult[93] = mult[29];
			temp_mult[94] = mult[30];
			temp_mult[95] = mult[31];
			temp_mult[96] = mult[32];
			temp_mult[97] = mult[33];
			temp_mult[98] = mult[34];
			temp_mult[99] = mult[35];
			temp_mult[100] =mult[36];
			temp_mult[101] =mult[37];
			temp_mult[102] =mult[38];
			temp_mult[103] =mult[39];
			temp_mult[104] =mult[40];
			temp_mult[105] =mult[41];
			temp_mult[106] =mult[42];
			temp_mult[107] =mult[43];
			temp_mult[108] =mult[44];
			temp_mult[109] =mult[45];
			temp_mult[110] =mult[46];
			temp_mult[111] =mult[47];
			temp_mult[112] =mult[48];
			temp_mult[113] =mult[49];
			temp_mult[114] =mult[50];
			temp_mult[115] =mult[51];
			temp_mult[116] =mult[52];
			temp_mult[117] =mult[53];
			temp_mult[118] =mult[54];
			temp_mult[119] =mult[55];
			temp_mult[120] =mult[56];
			temp_mult[121] =mult[57];
			temp_mult[122] =mult[58];
			temp_mult[123] =mult[59];
			temp_mult[124] =mult[60];
			temp_mult[125] =mult[61];
			temp_mult[126] =mult[62];
			temp_mult[127] =mult[63];
		end
		5'd3: begin
			b[0]  = d1_input_r[128];
			b[1]  = d1_input_r[129];
			b[2]  = d1_input_r[130];
			b[3]  = d1_input_r[131];
			b[4]  = d1_input_r[132];
			b[5]  = d1_input_r[133];
			b[6]  = d1_input_r[134];
			b[7]  = d1_input_r[135];
			b[8]  = d1_input_r[136];
			b[9]  = d1_input_r[137];
			b[10] = d1_input_r[138];
			b[11] = d1_input_r[139];
			b[12] = d1_input_r[140];
			b[13] = d1_input_r[141];
			b[14] = d1_input_r[142];
			b[15] = d1_input_r[143];
			b[16] = d1_input_r[144];
			b[17] = d1_input_r[145];
			b[18] = d1_input_r[146];
			b[19] = d1_input_r[147];
			b[20] = d1_input_r[148];
			b[21] = d1_input_r[149];
			b[22] = d1_input_r[150];
			b[23] = d1_input_r[151];
			b[24] = d1_input_r[152];
			b[25] = d1_input_r[153];
			b[26] = d1_input_r[154];
			b[27] = d1_input_r[155];
			b[28] = d1_input_r[156];
			b[29] = d1_input_r[157];
			b[30] = d1_input_r[158];
			b[31] = d1_input_r[159];
			b[32] = d1_input_r[160];
			b[33] = d1_input_r[161];
			b[34] = d1_input_r[162];
			b[35] = d1_input_r[163];
			b[36] = d1_input_r[164];
			b[37] = d1_input_r[165];
			b[38] = d1_input_r[166];
			b[39] = d1_input_r[167];
			b[40] = d1_input_r[168];
			b[41] = d1_input_r[169];
			b[42] = d1_input_r[170];
			b[43] = d1_input_r[171];
			b[44] = d1_input_r[172];
			b[45] = d1_input_r[173];
			b[46] = d1_input_r[174];
			b[47] = d1_input_r[175];
			b[48] = d1_input_r[176];
			b[49] = d1_input_r[177];
			b[50] = d1_input_r[178];
			b[51] = d1_input_r[179];
			b[52] = d1_input_r[180];
			b[53] = d1_input_r[181];
			b[54] = d1_input_r[182];
			b[55] = d1_input_r[183];
			b[56] = d1_input_r[184];
			b[57] = d1_input_r[185];
			b[58] = d1_input_r[186];
			b[59] = d1_input_r[187];
			b[60] = d1_input_r[188];
			b[61] = d1_input_r[189];
			b[62] = d1_input_r[190];
			b[63] = d1_input_r[191];
			a[0]  = 16'd1024 ;
			a[1]  = 16'd1619 ;
			a[2]  = 16'd1585 ;
			a[3]  = 16'd33496;
			a[4]  = 16'd34669;
			a[5]  = 16'd35444;
			a[6]  = 16'd34470;
			a[7]  = 16'd33334;
			a[8]  = 16'd2565 ;
			a[9]  = 16'd33420;
			a[10] = 16'd35502;
			a[11] = 16'd33781;
			a[12] = 16'd2085 ;
			a[13] = 16'd328  ;
			a[14] = 16'd32903;
			a[15] = 16'd33928;
			a[16] = 16'd34128;
			a[17] = 16'd34319;
			a[18] = 16'd33171;
			a[19] = 16'd34067;
			a[20] = 16'd381  ;
			a[21] = 16'd1803 ;
			a[22] = 16'd110  ;
			a[23] = 16'd33524;
			a[24] = 16'd33441;
			a[25] = 16'd1502 ;
			a[26] = 16'd1843 ;
			a[27] = 16'd33835;
			a[28] = 16'd1056 ;
			a[29] = 16'd573  ;
			a[30] = 16'd33310;
			a[31] = 16'd34185;
			a[32] = 16'd378  ;
			a[33] = 16'd32980;
			a[34] = 16'd318  ;
			a[35] = 16'd34115;
			a[36] = 16'd740  ;
			a[37] = 16'd33599;
			a[38] = 16'd34725;
			a[39] = 16'd555  ;
			a[40] = 16'd33489;
			a[41] = 16'd32988;
			a[42] = 16'd136  ;
			a[43] = 16'd33689;
			a[44] = 16'd32816;
			a[45] = 16'd1937 ;
			a[46] = 16'd33731;
			a[47] = 16'd1016 ;
			a[48] = 16'd1585 ;
			a[49] = 16'd462  ;
			a[50] = 16'd33246;
			a[51] = 16'd659  ;
			a[52] = 16'd35100;
			a[53] = 16'd33522;
			a[54] = 16'd781  ;
			a[55] = 16'd630  ;
			a[56] = 16'd32788;
			a[57] = 16'd33054;
			a[58] = 16'd2849 ;
			a[59] = 16'd2577 ;
			a[60] = 16'd33140;
			a[61] = 16'd1847 ;
			a[62] = 16'd33543;
			a[63] = 16'd1058 ;
			temp_mult[128] =mult[0] ;
			temp_mult[129] =mult[1] ;
			temp_mult[130] =mult[2] ;
			temp_mult[131] =mult[3] ;
			temp_mult[132] =mult[4] ;
			temp_mult[133] =mult[5] ;
			temp_mult[134] =mult[6] ;
			temp_mult[135] =mult[7] ;
			temp_mult[136] =mult[8] ;
			temp_mult[137] =mult[9] ;
			temp_mult[138] =mult[10];
			temp_mult[139] =mult[11];
			temp_mult[140] =mult[12];
			temp_mult[141] =mult[13];
			temp_mult[142] =mult[14];
			temp_mult[143] =mult[15];
			temp_mult[144] =mult[16];
			temp_mult[145] =mult[17];
			temp_mult[146] =mult[18];
			temp_mult[147] =mult[19];
			temp_mult[148] =mult[20];
			temp_mult[149] =mult[21];
			temp_mult[150] =mult[22];
			temp_mult[151] =mult[23];
			temp_mult[152] =mult[24];
			temp_mult[153] =mult[25];
			temp_mult[154] =mult[26];
			temp_mult[155] =mult[27];
			temp_mult[156] =mult[28];
			temp_mult[157] =mult[29];
			temp_mult[158] =mult[30];
			temp_mult[159] =mult[31];
			temp_mult[160] =mult[32];
			temp_mult[161] =mult[33];
			temp_mult[162] =mult[34];
			temp_mult[163] =mult[35];
			temp_mult[164] =mult[36];
			temp_mult[165] =mult[37];
			temp_mult[166] =mult[38];
			temp_mult[167] =mult[39];
			temp_mult[168] =mult[40];
			temp_mult[169] =mult[41];
			temp_mult[170] =mult[42];
			temp_mult[171] =mult[43];
			temp_mult[172] =mult[44];
			temp_mult[173] =mult[45];
			temp_mult[174] =mult[46];
			temp_mult[175] =mult[47];
			temp_mult[176] =mult[48];
			temp_mult[177] =mult[49];
			temp_mult[178] =mult[50];
			temp_mult[179] =mult[51];
			temp_mult[180] =mult[52];
			temp_mult[181] =mult[53];
			temp_mult[182] =mult[54];
			temp_mult[183] =mult[55];
			temp_mult[184] =mult[56];
			temp_mult[185] =mult[57];
			temp_mult[186] =mult[58];
			temp_mult[187] =mult[59];
			temp_mult[188] =mult[60];
			temp_mult[189] =mult[61];
			temp_mult[190] =mult[62];
			temp_mult[191] =mult[63];
		end
		5'd4: begin
			b[0]  = d1_input_r[192];
			b[1]  = d1_input_r[193];
			b[2]  = d1_input_r[194];
			b[3]  = d1_input_r[195];
			b[4]  = d1_input_r[196];
			b[5]  = d1_input_r[197];
			b[6]  = d1_input_r[198];
			b[7]  = d1_input_r[199];
			b[8]  = d1_input_r[200];
			b[9]  = d1_input_r[201];
			b[10] = d1_input_r[202];
			b[11] = d1_input_r[203];
			b[12] = d1_input_r[204];
			b[13] = d1_input_r[205];
			b[14] = d1_input_r[206];
			b[15] = d1_input_r[207];
			b[16] = d1_input_r[208];
			b[17] = d1_input_r[209];
			b[18] = d1_input_r[210];
			b[19] = d1_input_r[211];
			b[20] = d1_input_r[212];
			b[21] = d1_input_r[213];
			b[22] = d1_input_r[214];
			b[23] = d1_input_r[215];
			b[24] = d1_input_r[216];
			b[25] = d1_input_r[217];
			b[26] = d1_input_r[218];
			b[27] = d1_input_r[219];
			b[28] = d1_input_r[220];
			b[29] = d1_input_r[221];
			b[30] = d1_input_r[222];
			b[31] = d1_input_r[223];
			b[32] = d1_input_r[224];
			b[33] = d1_input_r[225];
			b[34] = d1_input_r[226];
			b[35] = d1_input_r[227];
			b[36] = d1_input_r[228];
			b[37] = d1_input_r[229];
			b[38] = d1_input_r[230];
			b[39] = d1_input_r[231];
			b[40] = d1_input_r[232];
			b[41] = d1_input_r[233];
			b[42] = d1_input_r[234];
			b[43] = d1_input_r[235];
			b[44] = d1_input_r[236];
			b[45] = d1_input_r[237];
			b[46] = d1_input_r[238];
			b[47] = d1_input_r[239];
			b[48] = d1_input_r[240];
			b[49] = d1_input_r[241];
			b[50] = d1_input_r[242];
			b[51] = d1_input_r[243];
			b[52] = d1_input_r[244];
			b[53] = d1_input_r[245];
			b[54] = d1_input_r[246];
			b[55] = d1_input_r[247];
			b[56] = d1_input_r[248];
			b[57] = d1_input_r[249];
			b[58] = d1_input_r[250];
			b[59] = d1_input_r[251];
			b[60] = d1_input_r[252];
			b[61] = d1_input_r[253];
			b[62] = d1_input_r[254];
			b[63] = d1_input_r[255];
			a[0]  = 16'd61   ;
			a[1]  = 16'd432  ;
			a[2]  = 16'd33782;
			a[3]  = 16'd33483;
			a[4]  = 16'd1453 ;
			a[5]  = 16'd1136 ;
			a[6]  = 16'd34849;
			a[7]  = 16'd2280 ;
			a[8]  = 16'd2566 ;
			a[9]  = 16'd34460;
			a[10] = 16'd34294;
			a[11] = 16'd1276 ;
			a[12] = 16'd1970 ;
			a[13] = 16'd34243;
			a[14] = 16'd1322 ;
			a[15] = 16'd34864;
			a[16] = 16'd33303;
			a[17] = 16'd407  ;
			a[18] = 16'd1732 ;
			a[19] = 16'd340  ;
			a[20] = 16'd1022 ;
			a[21] = 16'd34272;
			a[22] = 16'd33965;
			a[23] = 16'd1057 ;
			a[24] = 16'd215  ;
			a[25] = 16'd1738 ;
			a[26] = 16'd1293 ;
			a[27] = 16'd3146 ;
			a[28] = 16'd1060 ;
			a[29] = 16'd1543 ;
			a[30] = 16'd296  ;
			a[31] = 16'd33327;
			a[32] = 16'd34496;
			a[33] = 16'd33170;
			a[34] = 16'd507  ;
			a[35] = 16'd2815 ;
			a[36] = 16'd33973;
			a[37] = 16'd33730;
			a[38] = 16'd33450;
			a[39] = 16'd687  ;
			a[40] = 16'd2561 ;
			a[41] = 16'd34430;
			a[42] = 16'd802  ;
			a[43] = 16'd34961;
			a[44] = 16'd1664 ;
			a[45] = 16'd1431 ;
			a[46] = 16'd799  ;
			a[47] = 16'd34597;
			a[48] = 16'd35550;
			a[49] = 16'd831  ;
			a[50] = 16'd717  ;
			a[51] = 16'd33328;
			a[52] = 16'd35745;
			a[53] = 16'd33702;
			a[54] = 16'd632  ;
			a[55] = 16'd34382;
			a[56] = 16'd520  ;
			a[57] = 16'd1811 ;
			a[58] = 16'd33937;
			a[59] = 16'd2222 ;
			a[60] = 16'd1776 ;
			a[61] = 16'd862  ;
			a[62] = 16'd34076;
			a[63] = 16'd2403 ;
			temp_mult[192] =mult[0] ;
			temp_mult[193] =mult[1] ;
			temp_mult[194] =mult[2] ;
			temp_mult[195] =mult[3] ;
			temp_mult[196] =mult[4] ;
			temp_mult[197] =mult[5] ;
			temp_mult[198] =mult[6] ;
			temp_mult[199] =mult[7] ;
			temp_mult[200] =mult[8] ;
			temp_mult[201] =mult[9] ;
			temp_mult[202] =mult[10];
			temp_mult[203] =mult[11];
			temp_mult[204] =mult[12];
			temp_mult[205] =mult[13];
			temp_mult[206] =mult[14];
			temp_mult[207] =mult[15];
			temp_mult[208] =mult[16];
			temp_mult[209] =mult[17];
			temp_mult[210] =mult[18];
			temp_mult[211] =mult[19];
			temp_mult[212] =mult[20];
			temp_mult[213] =mult[21];
			temp_mult[214] =mult[22];
			temp_mult[215] =mult[23];
			temp_mult[216] =mult[24];
			temp_mult[217] =mult[25];
			temp_mult[218] =mult[26];
			temp_mult[219] =mult[27];
			temp_mult[220] =mult[28];
			temp_mult[221] =mult[29];
			temp_mult[222] =mult[30];
			temp_mult[223] =mult[31];
			temp_mult[224] =mult[32];
			temp_mult[225] =mult[33];
			temp_mult[226] =mult[34];
			temp_mult[227] =mult[35];
			temp_mult[228] =mult[36];
			temp_mult[229] =mult[37];
			temp_mult[230] =mult[38];
			temp_mult[231] =mult[39];
			temp_mult[232] =mult[40];
			temp_mult[233] =mult[41];
			temp_mult[234] =mult[42];
			temp_mult[235] =mult[43];
			temp_mult[236] =mult[44];
			temp_mult[237] =mult[45];
			temp_mult[238] =mult[46];
			temp_mult[239] =mult[47];
			temp_mult[240] =mult[48];
			temp_mult[241] =mult[49];
			temp_mult[242] =mult[50];
			temp_mult[243] =mult[51];
			temp_mult[244] =mult[52];
			temp_mult[245] =mult[53];
			temp_mult[246] =mult[54];
			temp_mult[247] =mult[55];
			temp_mult[248] =mult[56];
			temp_mult[249] =mult[57];
			temp_mult[250] =mult[58];
			temp_mult[251] =mult[59];
			temp_mult[252] =mult[60];
			temp_mult[253] =mult[61];
			temp_mult[254] =mult[62];
			temp_mult[255] =mult[63];
		end
		5'd5: begin
			b[0]  =  d1_input_r[0];
			b[1]  =  d1_input_r[1];
			b[2]  =  d1_input_r[2];
			b[3]  =  d1_input_r[3];
			b[4]  =  d1_input_r[4];
			b[5]  =  d1_input_r[5];
			b[6]  =  d1_input_r[6];
			b[7]  =  d1_input_r[7];
			b[8]  =  d1_input_r[8];
			b[9]  =  d1_input_r[9];
			b[10] =  d1_input_r[10];
			b[11] =  d1_input_r[11];
			b[12] =  d1_input_r[12];
			b[13] =  d1_input_r[13];
			b[14] =  d1_input_r[14];
			b[15] =  d1_input_r[15];
			b[16] =  d1_input_r[16];
			b[17] =  d1_input_r[17];
			b[18] =  d1_input_r[18];
			b[19] =  d1_input_r[19];
			b[20] =  d1_input_r[20];
			b[21] =  d1_input_r[21];
			b[22] =  d1_input_r[22];
			b[23] =  d1_input_r[23];
			b[24] =  d1_input_r[24];
			b[25] =  d1_input_r[25];
			b[26] =  d1_input_r[26];
			b[27] =  d1_input_r[27];
			b[28] =  d1_input_r[28];
			b[29] =  d1_input_r[29];
			b[30] =  d1_input_r[30];
			b[31] =  d1_input_r[31];
			b[32] =  d1_input_r[32];
			b[33] =  d1_input_r[33];
			b[34] =  d1_input_r[34];
			b[35] =  d1_input_r[35];
			b[36] =  d1_input_r[36];
			b[37] =  d1_input_r[37];
			b[38] =  d1_input_r[38];
			b[39] =  d1_input_r[39];
			b[40] =  d1_input_r[40];
			b[41] =  d1_input_r[41];
			b[42] =  d1_input_r[42];
			b[43] =  d1_input_r[43];
			b[44] =  d1_input_r[44];
			b[45] =  d1_input_r[45];
			b[46] =  d1_input_r[46];
			b[47] =  d1_input_r[47];
			b[48] =  d1_input_r[48];
			b[49] =  d1_input_r[49];
			b[50] =  d1_input_r[50];
			b[51] =  d1_input_r[51];
			b[52] =  d1_input_r[52];
			b[53] =  d1_input_r[53];
			b[54] =  d1_input_r[54];
			b[55] =  d1_input_r[55];
			b[56] =  d1_input_r[56];
			b[57] =  d1_input_r[57];
			b[58] =  d1_input_r[58];
			b[59] =  d1_input_r[59];
			b[60] =  d1_input_r[60];
			b[61] =  d1_input_r[61];
			b[62] =  d1_input_r[62];
			b[63] =  d1_input_r[63];
			a[0]  =16'd1741 ;
			a[1]  =16'd580  ;
			a[2]  =16'd644  ;
			a[3]  =16'd33412;
			a[4]  =16'd33545;
			a[5]  =16'd35146;
			a[6]  =16'd1832 ;
			a[7]  =16'd1903 ;
			a[8]  =16'd1961 ;
			a[9]  =16'd34914;
			a[10] =16'd2360 ;
			a[11] =16'd907  ;
			a[12] =16'd32869;
			a[13] =16'd33679;
			a[14] =16'd32944;
			a[15] =16'd600  ;
			a[16] =16'd1603 ;
			a[17] =16'd33544;
			a[18] =16'd35058;
			a[19] =16'd32895;
			a[20] =16'd33413;
			a[21] =16'd35193;
			a[22] =16'd858  ;
			a[23] =16'd1606 ;
			a[24] =16'd1359 ;
			a[25] =16'd359  ;
			a[26] =16'd1545 ;
			a[27] =16'd33911;
			a[28] =16'd132  ;
			a[29] =16'd35108;
			a[30] =16'd34614;
			a[31] =16'd33613;
			a[32] =16'd33508;
			a[33] =16'd1699 ;
			a[34] =16'd34507;
			a[35] =16'd2576 ;
			a[36] =16'd994  ;
			a[37] =16'd178  ;
			a[38] =16'd32786;
			a[39] =16'd33136;
			a[40] =16'd2550 ;
			a[41] =16'd34846;
			a[42] =16'd33587;
			a[43] =16'd34555;
			a[44] =16'd35646;
			a[45] =16'd34822;
			a[46] =16'd866  ;
			a[47] =16'd33467;
			a[48] =16'd1925 ;
			a[49] =16'd532  ;
			a[50] =16'd1213 ;
			a[51] =16'd1065 ;
			a[52] =16'd34078;
			a[53] =16'd33242;
			a[54] =16'd1949 ;
			a[55] =16'd33600;
			a[56] =16'd915  ;
			a[57] =16'd1177 ;
			a[58] =16'd34051;
			a[59] =16'd1066 ;
			a[60] =16'd1121 ;
			a[61] =16'd33143;
			a[62] =16'd34049;
			a[63] =16'd1024 ;
			temp_mult[256] =mult[0] ;
			temp_mult[257] =mult[1] ;
			temp_mult[258] =mult[2] ;
			temp_mult[259] =mult[3] ;
			temp_mult[260] =mult[4] ;
			temp_mult[261] =mult[5] ;
			temp_mult[262] =mult[6] ;
			temp_mult[263] =mult[7] ;
			temp_mult[264] =mult[8] ;
			temp_mult[265] =mult[9] ;
			temp_mult[266] =mult[10];
			temp_mult[267] =mult[11];
			temp_mult[268] =mult[12];
			temp_mult[269] =mult[13];
			temp_mult[270] =mult[14];
			temp_mult[271] =mult[15];
			temp_mult[272] =mult[16];
			temp_mult[273] =mult[17];
			temp_mult[274] =mult[18];
			temp_mult[275] =mult[19];
			temp_mult[276] =mult[20];
			temp_mult[277] =mult[21];
			temp_mult[278] =mult[22];
			temp_mult[279] =mult[23];
			temp_mult[280] =mult[24];
			temp_mult[281] =mult[25];
			temp_mult[282] =mult[26];
			temp_mult[283] =mult[27];
			temp_mult[284] =mult[28];
			temp_mult[285] =mult[29];
			temp_mult[286] =mult[30];
			temp_mult[287] =mult[31];
			temp_mult[288] =mult[32];
			temp_mult[289] =mult[33];
			temp_mult[290] =mult[34];
			temp_mult[291] =mult[35];
			temp_mult[292] =mult[36];
			temp_mult[293] =mult[37];
			temp_mult[294] =mult[38];
			temp_mult[295] =mult[39];
			temp_mult[296] =mult[40];
			temp_mult[297] =mult[41];
			temp_mult[298] =mult[42];
			temp_mult[299] =mult[43];
			temp_mult[300] =mult[44];
			temp_mult[301] =mult[45];
			temp_mult[302] =mult[46];
			temp_mult[303] =mult[47];
			temp_mult[304] =mult[48];
			temp_mult[305] =mult[49];
			temp_mult[306] =mult[50];
			temp_mult[307] =mult[51];
			temp_mult[308] =mult[52];
			temp_mult[309] =mult[53];
			temp_mult[310] =mult[54];
			temp_mult[311] =mult[55];
			temp_mult[312] =mult[56];
			temp_mult[313] =mult[57];
			temp_mult[314] =mult[58];
			temp_mult[315] =mult[59];
			temp_mult[316] =mult[60];
			temp_mult[317] =mult[61];
			temp_mult[318] =mult[62];
			temp_mult[319] =mult[63];
		end
		5'd6: begin
			b[0]  = d1_input_r[64];
			b[1]  = d1_input_r[65];
			b[2]  = d1_input_r[66];
			b[3]  = d1_input_r[67];
			b[4]  = d1_input_r[68];
			b[5]  = d1_input_r[69];
			b[6]  = d1_input_r[70];
			b[7]  = d1_input_r[71];
			b[8]  = d1_input_r[72];
			b[9]  = d1_input_r[73];
			b[10] = d1_input_r[74];
			b[11] = d1_input_r[75];
			b[12] = d1_input_r[76];
			b[13] = d1_input_r[77];
			b[14] = d1_input_r[78];
			b[15] = d1_input_r[79];
			b[16] = d1_input_r[80];
			b[17] = d1_input_r[81];
			b[18] = d1_input_r[82];
			b[19] = d1_input_r[83];
			b[20] = d1_input_r[84];
			b[21] = d1_input_r[85];
			b[22] = d1_input_r[86];
			b[23] = d1_input_r[87];
			b[24] = d1_input_r[88];
			b[25] = d1_input_r[89];
			b[26] = d1_input_r[90];
			b[27] = d1_input_r[91];
			b[28] = d1_input_r[92];
			b[29] = d1_input_r[93];
			b[30] = d1_input_r[94];
			b[31] = d1_input_r[95];
			b[32] = d1_input_r[96];
			b[33] = d1_input_r[97];
			b[34] = d1_input_r[98];
			b[35] = d1_input_r[99];
			b[36] = d1_input_r[100];
			b[37] = d1_input_r[101];
			b[38] = d1_input_r[102];
			b[39] = d1_input_r[103];
			b[40] = d1_input_r[104];
			b[41] = d1_input_r[105];
			b[42] = d1_input_r[106];
			b[43] = d1_input_r[107];
			b[44] = d1_input_r[108];
			b[45] = d1_input_r[109];
			b[46] = d1_input_r[110];
			b[47] = d1_input_r[111];
			b[48] = d1_input_r[112];
			b[49] = d1_input_r[113];
			b[50] = d1_input_r[114];
			b[51] = d1_input_r[115];
			b[52] = d1_input_r[116];
			b[53] = d1_input_r[117];
			b[54] = d1_input_r[118];
			b[55] = d1_input_r[119];
			b[56] = d1_input_r[120];
			b[57] = d1_input_r[121];
			b[58] = d1_input_r[122];
			b[59] = d1_input_r[123];
			b[60] = d1_input_r[124];
			b[61] = d1_input_r[125];
			b[62] = d1_input_r[126];
			b[63] = d1_input_r[127];
			a[0]  =16'd449  ;
			a[1]  =16'd34668;
			a[2]  =16'd175  ;
			a[3]  =16'd34370;
			a[4]  =16'd131  ;
			a[5]  =16'd34900;
			a[6]  =16'd169  ;
			a[7]  =16'd1022 ;
			a[8]  =16'd767  ;
			a[9]  =16'd35378;
			a[10] =16'd106  ;
			a[11] =16'd964  ;
			a[12] =16'd33114;
			a[13] =16'd407  ;
			a[14] =16'd1887 ;
			a[15] =16'd35161;
			a[16] =16'd34277;
			a[17] =16'd962  ;
			a[18] =16'd1023 ;
			a[19] =16'd35844;
			a[20] =16'd1524 ;
			a[21] =16'd3028 ;
			a[22] =16'd33678;
			a[23] =16'd33406;
			a[24] =16'd1591 ;
			a[25] =16'd1445 ;
			a[26] =16'd34257;
			a[27] =16'd33017;
			a[28] =16'd184  ;
			a[29] =16'd811  ;
			a[30] =16'd34839;
			a[31] =16'd2238 ;
			a[32] =16'd34491;
			a[33] =16'd579  ;
			a[34] =16'd1670 ;
			a[35] =16'd1554 ;
			a[36] =16'd34742;
			a[37] =16'd1031 ;
			a[38] =16'd1224 ;
			a[39] =16'd2158 ;
			a[40] =16'd1880 ;
			a[41] =16'd32913;
			a[42] =16'd33427;
			a[43] =16'd2340 ;
			a[44] =16'd34072;
			a[45] =16'd32983;
			a[46] =16'd34055;
			a[47] =16'd544  ;
			a[48] =16'd34468;
			a[49] =16'd2794 ;
			a[50] =16'd32841;
			a[51] =16'd33397;
			a[52] =16'd605  ;
			a[53] =16'd33916;
			a[54] =16'd33556;
			a[55] =16'd34927;
			a[56] =16'd580  ;
			a[57] =16'd1346 ;
			a[58] =16'd530  ;
			a[59] =16'd33930;
			a[60] =16'd1364 ;
			a[61] =16'd1351 ;
			a[62] =16'd2027 ;
			a[63] =16'd33636;
			temp_mult[320] = mult[0] ;
			temp_mult[321] = mult[1] ;
			temp_mult[322] = mult[2] ;
			temp_mult[323] = mult[3] ;
			temp_mult[324] = mult[4] ;
			temp_mult[325] = mult[5] ;
			temp_mult[326] = mult[6] ;
			temp_mult[327] = mult[7] ;
			temp_mult[328] = mult[8] ;
			temp_mult[329] = mult[9] ;
			temp_mult[330] = mult[10];
			temp_mult[331] = mult[11];
			temp_mult[332] = mult[12];
			temp_mult[333] = mult[13];
			temp_mult[334] = mult[14];
			temp_mult[335] = mult[15];
			temp_mult[336] = mult[16];
			temp_mult[337] = mult[17];
			temp_mult[338] = mult[18];
			temp_mult[339] = mult[19];
			temp_mult[340] = mult[20];
			temp_mult[341] = mult[21];
			temp_mult[342] = mult[22];
			temp_mult[343] = mult[23];
			temp_mult[344] = mult[24];
			temp_mult[345] = mult[25];
			temp_mult[346] = mult[26];
			temp_mult[347] = mult[27];
			temp_mult[348] = mult[28];
			temp_mult[349] = mult[29];
			temp_mult[350] = mult[30];
			temp_mult[351] = mult[31];
			temp_mult[352] = mult[32];
			temp_mult[353] = mult[33];
			temp_mult[354] = mult[34];
			temp_mult[355] = mult[35];
			temp_mult[356] = mult[36];
			temp_mult[357] = mult[37];
			temp_mult[358] = mult[38];
			temp_mult[359] = mult[39];
			temp_mult[360] = mult[40];
			temp_mult[361] = mult[41];
			temp_mult[362] = mult[42];
			temp_mult[363] = mult[43];
			temp_mult[364] = mult[44];
			temp_mult[365] = mult[45];
			temp_mult[366] = mult[46];
			temp_mult[367] = mult[47];
			temp_mult[368] = mult[48];
			temp_mult[369] = mult[49];
			temp_mult[370] = mult[50];
			temp_mult[371] = mult[51];
			temp_mult[372] = mult[52];
			temp_mult[373] = mult[53];
			temp_mult[374] = mult[54];
			temp_mult[375] = mult[55];
			temp_mult[376] = mult[56];
			temp_mult[377] = mult[57];
			temp_mult[378] = mult[58];
			temp_mult[379] = mult[59];
			temp_mult[380] = mult[60];
			temp_mult[381] = mult[61];
			temp_mult[382] = mult[62];
			temp_mult[383] = mult[63];
		end
		5'd7: begin
			b[0]  = d1_input_r[128];
			b[1]  = d1_input_r[129];
			b[2]  = d1_input_r[130];
			b[3]  = d1_input_r[131];
			b[4]  = d1_input_r[132];
			b[5]  = d1_input_r[133];
			b[6]  = d1_input_r[134];
			b[7]  = d1_input_r[135];
			b[8]  = d1_input_r[136];
			b[9]  = d1_input_r[137];
			b[10] = d1_input_r[138];
			b[11] = d1_input_r[139];
			b[12] = d1_input_r[140];
			b[13] = d1_input_r[141];
			b[14] = d1_input_r[142];
			b[15] = d1_input_r[143];
			b[16] = d1_input_r[144];
			b[17] = d1_input_r[145];
			b[18] = d1_input_r[146];
			b[19] = d1_input_r[147];
			b[20] = d1_input_r[148];
			b[21] = d1_input_r[149];
			b[22] = d1_input_r[150];
			b[23] = d1_input_r[151];
			b[24] = d1_input_r[152];
			b[25] = d1_input_r[153];
			b[26] = d1_input_r[154];
			b[27] = d1_input_r[155];
			b[28] = d1_input_r[156];
			b[29] = d1_input_r[157];
			b[30] = d1_input_r[158];
			b[31] = d1_input_r[159];
			b[32] = d1_input_r[160];
			b[33] = d1_input_r[161];
			b[34] = d1_input_r[162];
			b[35] = d1_input_r[163];
			b[36] = d1_input_r[164];
			b[37] = d1_input_r[165];
			b[38] = d1_input_r[166];
			b[39] = d1_input_r[167];
			b[40] = d1_input_r[168];
			b[41] = d1_input_r[169];
			b[42] = d1_input_r[170];
			b[43] = d1_input_r[171];
			b[44] = d1_input_r[172];
			b[45] = d1_input_r[173];
			b[46] = d1_input_r[174];
			b[47] = d1_input_r[175];
			b[48] = d1_input_r[176];
			b[49] = d1_input_r[177];
			b[50] = d1_input_r[178];
			b[51] = d1_input_r[179];
			b[52] = d1_input_r[180];
			b[53] = d1_input_r[181];
			b[54] = d1_input_r[182];
			b[55] = d1_input_r[183];
			b[56] = d1_input_r[184];
			b[57] = d1_input_r[185];
			b[58] = d1_input_r[186];
			b[59] = d1_input_r[187];
			b[60] = d1_input_r[188];
			b[61] = d1_input_r[189];
			b[62] = d1_input_r[190];
			b[63] = d1_input_r[191];
			a[0]  =16'd420  ;
			a[1]  =16'd35008;
			a[2]  =16'd34166;
			a[3]  =16'd33450;
			a[4]  =16'd34803;
			a[5]  =16'd35081;
			a[6]  =16'd35312;
			a[7]  =16'd3088 ;
			a[8]  =16'd2911 ;
			a[9]  =16'd1473 ;
			a[10] =16'd1851 ;
			a[11] =16'd752  ;
			a[12] =16'd33051;
			a[13] =16'd2588 ;
			a[14] =16'd9    ;
			a[15] =16'd919  ;
			a[16] =16'd82   ;
			a[17] =16'd1822 ;
			a[18] =16'd33799;
			a[19] =16'd35337;
			a[20] =16'd1641 ;
			a[21] =16'd34106;
			a[22] =16'd33158;
			a[23] =16'd534  ;
			a[24] =16'd1553 ;
			a[25] =16'd35250;
			a[26] =16'd552  ;
			a[27] =16'd1387 ;
			a[28] =16'd2896 ;
			a[29] =16'd33531;
			a[30] =16'd34582;
			a[31] =16'd590  ;
			a[32] =16'd34816;
			a[33] =16'd34292;
			a[34] =16'd90   ;
			a[35] =16'd1120 ;
			a[36] =16'd416  ;
			a[37] =16'd34664;
			a[38] =16'd543  ;
			a[39] =16'd2847 ;
			a[40] =16'd1904 ;
			a[41] =16'd34336;
			a[42] =16'd34073;
			a[43] =16'd33829;
			a[44] =16'd13   ;
			a[45] =16'd454  ;
			a[46] =16'd34606;
			a[47] =16'd32777;
			a[48] =16'd150  ;
			a[49] =16'd32839;
			a[50] =16'd1999 ;
			a[51] =16'd34879;
			a[52] =16'd63   ;
			a[53] =16'd33351;
			a[54] =16'd393  ;
			a[55] =16'd33995;
			a[56] =16'd895  ;
			a[57] =16'd1694 ;
			a[58] =16'd248  ;
			a[59] =16'd33020;
			a[60] =16'd32832;
			a[61] =16'd33787;
			a[62] =16'd35556;
			a[63] =16'd32810;
			temp_mult[384] = mult[0] ;
			temp_mult[385] = mult[1] ;
			temp_mult[386] = mult[2] ;
			temp_mult[387] = mult[3] ;
			temp_mult[388] = mult[4] ;
			temp_mult[389] = mult[5] ;
			temp_mult[390] = mult[6] ;
			temp_mult[391] = mult[7] ;
			temp_mult[392] = mult[8] ;
			temp_mult[393] = mult[9] ;
			temp_mult[394] = mult[10];
			temp_mult[395] = mult[11];
			temp_mult[396] = mult[12];
			temp_mult[397] = mult[13];
			temp_mult[398] = mult[14];
			temp_mult[399] = mult[15];
			temp_mult[400] = mult[16];
			temp_mult[401] = mult[17];
			temp_mult[402] = mult[18];
			temp_mult[403] = mult[19];
			temp_mult[404] = mult[20];
			temp_mult[405] = mult[21];
			temp_mult[406] = mult[22];
			temp_mult[407] = mult[23];
			temp_mult[408] = mult[24];
			temp_mult[409] = mult[25];
			temp_mult[410] = mult[26];
			temp_mult[411] = mult[27];
			temp_mult[412] = mult[28];
			temp_mult[413] = mult[29];
			temp_mult[414] = mult[30];
			temp_mult[415] = mult[31];
			temp_mult[416] = mult[32];
			temp_mult[417] = mult[33];
			temp_mult[418] = mult[34];
			temp_mult[419] = mult[35];
			temp_mult[420] = mult[36];
			temp_mult[421] = mult[37];
			temp_mult[422] = mult[38];
			temp_mult[423] = mult[39];
			temp_mult[424] = mult[40];
			temp_mult[425] = mult[41];
			temp_mult[426] = mult[42];
			temp_mult[427] = mult[43];
			temp_mult[428] = mult[44];
			temp_mult[429] = mult[45];
			temp_mult[430] = mult[46];
			temp_mult[431] = mult[47];
			temp_mult[432] = mult[48];
			temp_mult[433] = mult[49];
			temp_mult[434] = mult[50];
			temp_mult[435] = mult[51];
			temp_mult[436] = mult[52];
			temp_mult[437] = mult[53];
			temp_mult[438] = mult[54];
			temp_mult[439] = mult[55];
			temp_mult[440] = mult[56];
			temp_mult[441] = mult[57];
			temp_mult[442] = mult[58];
			temp_mult[443] = mult[59];
			temp_mult[444] = mult[60];
			temp_mult[445] = mult[61];
			temp_mult[446] = mult[62];
			temp_mult[447] = mult[63];
		end
		5'd8: begin
			b[0]  = d1_input_r[192];
			b[1]  = d1_input_r[193];
			b[2]  = d1_input_r[194];
			b[3]  = d1_input_r[195];
			b[4]  = d1_input_r[196];
			b[5]  = d1_input_r[197];
			b[6]  = d1_input_r[198];
			b[7]  = d1_input_r[199];
			b[8]  = d1_input_r[200];
			b[9]  = d1_input_r[201];
			b[10] = d1_input_r[202];
			b[11] = d1_input_r[203];
			b[12] = d1_input_r[204];
			b[13] = d1_input_r[205];
			b[14] = d1_input_r[206];
			b[15] = d1_input_r[207];
			b[16] = d1_input_r[208];
			b[17] = d1_input_r[209];
			b[18] = d1_input_r[210];
			b[19] = d1_input_r[211];
			b[20] = d1_input_r[212];
			b[21] = d1_input_r[213];
			b[22] = d1_input_r[214];
			b[23] = d1_input_r[215];
			b[24] = d1_input_r[216];
			b[25] = d1_input_r[217];
			b[26] = d1_input_r[218];
			b[27] = d1_input_r[219];
			b[28] = d1_input_r[220];
			b[29] = d1_input_r[221];
			b[30] = d1_input_r[222];
			b[31] = d1_input_r[223];
			b[32] = d1_input_r[224];
			b[33] = d1_input_r[225];
			b[34] = d1_input_r[226];
			b[35] = d1_input_r[227];
			b[36] = d1_input_r[228];
			b[37] = d1_input_r[229];
			b[38] = d1_input_r[230];
			b[39] = d1_input_r[231];
			b[40] = d1_input_r[232];
			b[41] = d1_input_r[233];
			b[42] = d1_input_r[234];
			b[43] = d1_input_r[235];
			b[44] = d1_input_r[236];
			b[45] = d1_input_r[237];
			b[46] = d1_input_r[238];
			b[47] = d1_input_r[239];
			b[48] = d1_input_r[240];
			b[49] = d1_input_r[241];
			b[50] = d1_input_r[242];
			b[51] = d1_input_r[243];
			b[52] = d1_input_r[244];
			b[53] = d1_input_r[245];
			b[54] = d1_input_r[246];
			b[55] = d1_input_r[247];
			b[56] = d1_input_r[248];
			b[57] = d1_input_r[249];
			b[58] = d1_input_r[250];
			b[59] = d1_input_r[251];
			b[60] = d1_input_r[252];
			b[61] = d1_input_r[253];
			b[62] = d1_input_r[254];
			b[63] = d1_input_r[255];
			a[0]  =16'd34013;
			a[1]  =16'd32872;
			a[2]  =16'd34942;
			a[3]  =16'd2430 ;
			a[4]  =16'd3005 ;
			a[5]  =16'd1292 ;
			a[6]  =16'd480  ;
			a[7]  =16'd33888;
			a[8]  =16'd149  ;
			a[9]  =16'd33879;
			a[10] =16'd776  ;
			a[11] =16'd34760;
			a[12] =16'd545  ;
			a[13] =16'd33914;
			a[14] =16'd34264;
			a[15] =16'd32956;
			a[16] =16'd35715;
			a[17] =16'd33075;
			a[18] =16'd1946 ;
			a[19] =16'd2275 ;
			a[20] =16'd239  ;
			a[21] =16'd35785;
			a[22] =16'd33729;
			a[23] =16'd691  ;
			a[24] =16'd1719 ;
			a[25] =16'd34842;
			a[26] =16'd33631;
			a[27] =16'd2998 ;
			a[28] =16'd73   ;
			a[29] =16'd1222 ;
			a[30] =16'd35619;
			a[31] =16'd1577 ;
			a[32] =16'd327  ;
			a[33] =16'd921  ;
			a[34] =16'd33839;
			a[35] =16'd2244 ;
			a[36] =16'd33637;
			a[37] =16'd33625;
			a[38] =16'd1644 ;
			a[39] =16'd33886;
			a[40] =16'd34508;
			a[41] =16'd33641;
			a[42] =16'd678  ;
			a[43] =16'd1838 ;
			a[44] =16'd34908;
			a[45] =16'd2054 ;
			a[46] =16'd802  ;
			a[47] =16'd34375;
			a[48] =16'd1084 ;
			a[49] =16'd1963 ;
			a[50] =16'd34540;
			a[51] =16'd1779 ;
			a[52] =16'd33956;
			a[53] =16'd33525;
			a[54] =16'd208  ;
			a[55] =16'd32888;
			a[56] =16'd1170 ;
			a[57] =16'd35266;
			a[58] =16'd620  ;
			a[59] =16'd344  ;
			a[60] =16'd1267 ;
			a[61] =16'd1764 ;
			a[62] =16'd33316;
			a[63] =16'd34   ;
			temp_mult[448] = mult[0] ;
			temp_mult[449] = mult[1] ;
			temp_mult[450] = mult[2] ;
			temp_mult[451] = mult[3] ;
			temp_mult[452] = mult[4] ;
			temp_mult[453] = mult[5] ;
			temp_mult[454] = mult[6] ;
			temp_mult[455] = mult[7] ;
			temp_mult[456] = mult[8] ;
			temp_mult[457] = mult[9] ;
			temp_mult[458] = mult[10];
			temp_mult[459] = mult[11];
			temp_mult[460] = mult[12];
			temp_mult[461] = mult[13];
			temp_mult[462] = mult[14];
			temp_mult[463] = mult[15];
			temp_mult[464] = mult[16];
			temp_mult[465] = mult[17];
			temp_mult[466] = mult[18];
			temp_mult[467] = mult[19];
			temp_mult[468] = mult[20];
			temp_mult[469] = mult[21];
			temp_mult[470] = mult[22];
			temp_mult[471] = mult[23];
			temp_mult[472] = mult[24];
			temp_mult[473] = mult[25];
			temp_mult[474] = mult[26];
			temp_mult[475] = mult[27];
			temp_mult[476] = mult[28];
			temp_mult[477] = mult[29];
			temp_mult[478] = mult[30];
			temp_mult[479] = mult[31];
			temp_mult[480] = mult[32];
			temp_mult[481] = mult[33];
			temp_mult[482] = mult[34];
			temp_mult[483] = mult[35];
			temp_mult[484] = mult[36];
			temp_mult[485] = mult[37];
			temp_mult[486] = mult[38];
			temp_mult[487] = mult[39];
			temp_mult[488] = mult[40];
			temp_mult[489] = mult[41];
			temp_mult[490] = mult[42];
			temp_mult[491] = mult[43];
			temp_mult[492] = mult[44];
			temp_mult[493] = mult[45];
			temp_mult[494] = mult[46];
			temp_mult[495] = mult[47];
			temp_mult[496] = mult[48];
			temp_mult[497] = mult[49];
			temp_mult[498] = mult[50];
			temp_mult[499] = mult[51];
			temp_mult[500] = mult[52];
			temp_mult[501] = mult[53];
			temp_mult[502] = mult[54];
			temp_mult[503] = mult[55];
			temp_mult[504] = mult[56];
			temp_mult[505] = mult[57];
			temp_mult[506] = mult[58];
			temp_mult[507] = mult[59];
			temp_mult[508] = mult[60];
			temp_mult[509] = mult[61];
			temp_mult[510] = mult[62];
			temp_mult[511] = mult[63];
		end
		5'd9: begin
			b[0]  =  d1_input_r[0];
			b[1]  =  d1_input_r[1];
			b[2]  =  d1_input_r[2];
			b[3]  =  d1_input_r[3];
			b[4]  =  d1_input_r[4];
			b[5]  =  d1_input_r[5];
			b[6]  =  d1_input_r[6];
			b[7]  =  d1_input_r[7];
			b[8]  =  d1_input_r[8];
			b[9]  =  d1_input_r[9];
			b[10] =  d1_input_r[10];
			b[11] =  d1_input_r[11];
			b[12] =  d1_input_r[12];
			b[13] =  d1_input_r[13];
			b[14] =  d1_input_r[14];
			b[15] =  d1_input_r[15];
			b[16] =  d1_input_r[16];
			b[17] =  d1_input_r[17];
			b[18] =  d1_input_r[18];
			b[19] =  d1_input_r[19];
			b[20] =  d1_input_r[20];
			b[21] =  d1_input_r[21];
			b[22] =  d1_input_r[22];
			b[23] =  d1_input_r[23];
			b[24] =  d1_input_r[24];
			b[25] =  d1_input_r[25];
			b[26] =  d1_input_r[26];
			b[27] =  d1_input_r[27];
			b[28] =  d1_input_r[28];
			b[29] =  d1_input_r[29];
			b[30] =  d1_input_r[30];
			b[31] =  d1_input_r[31];
			b[32] =  d1_input_r[32];
			b[33] =  d1_input_r[33];
			b[34] =  d1_input_r[34];
			b[35] =  d1_input_r[35];
			b[36] =  d1_input_r[36];
			b[37] =  d1_input_r[37];
			b[38] =  d1_input_r[38];
			b[39] =  d1_input_r[39];
			b[40] =  d1_input_r[40];
			b[41] =  d1_input_r[41];
			b[42] =  d1_input_r[42];
			b[43] =  d1_input_r[43];
			b[44] =  d1_input_r[44];
			b[45] =  d1_input_r[45];
			b[46] =  d1_input_r[46];
			b[47] =  d1_input_r[47];
			b[48] =  d1_input_r[48];
			b[49] =  d1_input_r[49];
			b[50] =  d1_input_r[50];
			b[51] =  d1_input_r[51];
			b[52] =  d1_input_r[52];
			b[53] =  d1_input_r[53];
			b[54] =  d1_input_r[54];
			b[55] =  d1_input_r[55];
			b[56] =  d1_input_r[56];
			b[57] =  d1_input_r[57];
			b[58] =  d1_input_r[58];
			b[59] =  d1_input_r[59];
			b[60] =  d1_input_r[60];
			b[61] =  d1_input_r[61];
			b[62] =  d1_input_r[62];
			b[63] =  d1_input_r[63];
			a[0]  =16'd34854;
			a[1]  =16'd32894;
			a[2]  =16'd33087;
			a[3]  =16'd35780;
			a[4]  =16'd32938;
			a[5]  =16'd3115 ;
			a[6]  =16'd33788;
			a[7]  =16'd1665 ;
			a[8]  =16'd255  ;
			a[9]  =16'd33302;
			a[10] =16'd35635;
			a[11] =16'd1048 ;
			a[12] =16'd32993;
			a[13] =16'd33350;
			a[14] =16'd34291;
			a[15] =16'd34515;
			a[16] =16'd2179 ;
			a[17] =16'd150  ;
			a[18] =16'd2025 ;
			a[19] =16'd33532;
			a[20] =16'd33189;
			a[21] =16'd1410 ;
			a[22] =16'd548  ;
			a[23] =16'd36   ;
			a[24] =16'd33979;
			a[25] =16'd878  ;
			a[26] =16'd2624 ;
			a[27] =16'd964  ;
			a[28] =16'd1693 ;
			a[29] =16'd906  ;
			a[30] =16'd1792 ;
			a[31] =16'd35761;
			a[32] =16'd33414;
			a[33] =16'd1335 ;
			a[34] =16'd34930;
			a[35] =16'd34174;
			a[36] =16'd1260 ;
			a[37] =16'd33425;
			a[38] =16'd35336;
			a[39] =16'd1229 ;
			a[40] =16'd1304 ;
			a[41] =16'd196  ;
			a[42] =16'd506  ;
			a[43] =16'd35113;
			a[44] =16'd2856 ;
			a[45] =16'd1360 ;
			a[46] =16'd34558;
			a[47] =16'd34245;
			a[48] =16'd829  ;
			a[49] =16'd126  ;
			a[50] =16'd32871;
			a[51] =16'd118  ;
			a[52] =16'd33735;
			a[53] =16'd34828;
			a[54] =16'd33243;
			a[55] =16'd2425 ;
			a[56] =16'd35539;
			a[57] =16'd34095;
			a[58] =16'd33530;
			a[59] =16'd34354;
			a[60] =16'd33064;
			a[61] =16'd1119 ;
			a[62] =16'd34288;
			a[63] =16'd754  ;
			temp_mult[512] = mult[0] ;
			temp_mult[513] = mult[1] ;
			temp_mult[514] = mult[2] ;
			temp_mult[515] = mult[3] ;
			temp_mult[516] = mult[4] ;
			temp_mult[517] = mult[5] ;
			temp_mult[518] = mult[6] ;
			temp_mult[519] = mult[7] ;
			temp_mult[520] = mult[8] ;
			temp_mult[521] = mult[9] ;
			temp_mult[522] = mult[10];
			temp_mult[523] = mult[11];
			temp_mult[524] = mult[12];
			temp_mult[525] = mult[13];
			temp_mult[526] = mult[14];
			temp_mult[527] = mult[15];
			temp_mult[528] = mult[16];
			temp_mult[529] = mult[17];
			temp_mult[530] = mult[18];
			temp_mult[531] = mult[19];
			temp_mult[532] = mult[20];
			temp_mult[533] = mult[21];
			temp_mult[534] = mult[22];
			temp_mult[535] = mult[23];
			temp_mult[536] = mult[24];
			temp_mult[537] = mult[25];
			temp_mult[538] = mult[26];
			temp_mult[539] = mult[27];
			temp_mult[540] = mult[28];
			temp_mult[541] = mult[29];
			temp_mult[542] = mult[30];
			temp_mult[543] = mult[31];
			temp_mult[544] = mult[32];
			temp_mult[545] = mult[33];
			temp_mult[546] = mult[34];
			temp_mult[547] = mult[35];
			temp_mult[548] = mult[36];
			temp_mult[549] = mult[37];
			temp_mult[550] = mult[38];
			temp_mult[551] = mult[39];
			temp_mult[552] = mult[40];
			temp_mult[553] = mult[41];
			temp_mult[554] = mult[42];
			temp_mult[555] = mult[43];
			temp_mult[556] = mult[44];
			temp_mult[557] = mult[45];
			temp_mult[558] = mult[46];
			temp_mult[559] = mult[47];
			temp_mult[560] = mult[48];
			temp_mult[561] = mult[49];
			temp_mult[562] = mult[50];
			temp_mult[563] = mult[51];
			temp_mult[564] = mult[52];
			temp_mult[565] = mult[53];
			temp_mult[566] = mult[54];
			temp_mult[567] = mult[55];
			temp_mult[568] = mult[56];
			temp_mult[569] = mult[57];
			temp_mult[570] = mult[58];
			temp_mult[571] = mult[59];
			temp_mult[572] = mult[60];
			temp_mult[573] = mult[61];
			temp_mult[574] = mult[62];
			temp_mult[575] = mult[63];
		end
		5'd10: begin
			b[0]  = d1_input_r[64];
			b[1]  = d1_input_r[65];
			b[2]  = d1_input_r[66];
			b[3]  = d1_input_r[67];
			b[4]  = d1_input_r[68];
			b[5]  = d1_input_r[69];
			b[6]  = d1_input_r[70];
			b[7]  = d1_input_r[71];
			b[8]  = d1_input_r[72];
			b[9]  = d1_input_r[73];
			b[10] = d1_input_r[74];
			b[11] = d1_input_r[75];
			b[12] = d1_input_r[76];
			b[13] = d1_input_r[77];
			b[14] = d1_input_r[78];
			b[15] = d1_input_r[79];
			b[16] = d1_input_r[80];
			b[17] = d1_input_r[81];
			b[18] = d1_input_r[82];
			b[19] = d1_input_r[83];
			b[20] = d1_input_r[84];
			b[21] = d1_input_r[85];
			b[22] = d1_input_r[86];
			b[23] = d1_input_r[87];
			b[24] = d1_input_r[88];
			b[25] = d1_input_r[89];
			b[26] = d1_input_r[90];
			b[27] = d1_input_r[91];
			b[28] = d1_input_r[92];
			b[29] = d1_input_r[93];
			b[30] = d1_input_r[94];
			b[31] = d1_input_r[95];
			b[32] = d1_input_r[96];
			b[33] = d1_input_r[97];
			b[34] = d1_input_r[98];
			b[35] = d1_input_r[99];
			b[36] = d1_input_r[100];
			b[37] = d1_input_r[101];
			b[38] = d1_input_r[102];
			b[39] = d1_input_r[103];
			b[40] = d1_input_r[104];
			b[41] = d1_input_r[105];
			b[42] = d1_input_r[106];
			b[43] = d1_input_r[107];
			b[44] = d1_input_r[108];
			b[45] = d1_input_r[109];
			b[46] = d1_input_r[110];
			b[47] = d1_input_r[111];
			b[48] = d1_input_r[112];
			b[49] = d1_input_r[113];
			b[50] = d1_input_r[114];
			b[51] = d1_input_r[115];
			b[52] = d1_input_r[116];
			b[53] = d1_input_r[117];
			b[54] = d1_input_r[118];
			b[55] = d1_input_r[119];
			b[56] = d1_input_r[120];
			b[57] = d1_input_r[121];
			b[58] = d1_input_r[122];
			b[59] = d1_input_r[123];
			b[60] = d1_input_r[124];
			b[61] = d1_input_r[125];
			b[62] = d1_input_r[126];
			b[63] = d1_input_r[127];
			a[0]  =16'd33814;
			a[1]  =16'd33496;
			a[2]  =16'd1002 ;
			a[3]  =16'd35658;
			a[4]  =16'd34031;
			a[5]  =16'd2293 ;
			a[6]  =16'd1847 ;
			a[7]  =16'd34447;
			a[8]  =16'd34904;
			a[9]  =16'd1708 ;
			a[10] =16'd33147;
			a[11] =16'd814  ;
			a[12] =16'd2926 ;
			a[13] =16'd2192 ;
			a[14] =16'd689  ;
			a[15] =16'd33769;
			a[16] =16'd33866;
			a[17] =16'd34800;
			a[18] =16'd33957;
			a[19] =16'd2888 ;
			a[20] =16'd34461;
			a[21] =16'd35748;
			a[22] =16'd1750 ;
			a[23] =16'd32950;
			a[24] =16'd35135;
			a[25] =16'd600  ;
			a[26] =16'd1379 ;
			a[27] =16'd35741;
			a[28] =16'd34353;
			a[29] =16'd2396 ;
			a[30] =16'd859  ;
			a[31] =16'd34582;
			a[32] =16'd646  ;
			a[33] =16'd1326 ;
			a[34] =16'd35144;
			a[35] =16'd33240;
			a[36] =16'd33956;
			a[37] =16'd32832;
			a[38] =16'd34316;
			a[39] =16'd698  ;
			a[40] =16'd1393 ;
			a[41] =16'd1141 ;
			a[42] =16'd972  ;
			a[43] =16'd34911;
			a[44] =16'd32945;
			a[45] =16'd1092 ;
			a[46] =16'd33433;
			a[47] =16'd33893;
			a[48] =16'd32849;
			a[49] =16'd35215;
			a[50] =16'd34464;
			a[51] =16'd1878 ;
			a[52] =16'd33327;
			a[53] =16'd722  ;
			a[54] =16'd35433;
			a[55] =16'd791  ;
			a[56] =16'd100  ;
			a[57] =16'd34389;
			a[58] =16'd33590;
			a[59] =16'd35287;
			a[60] =16'd35240;
			a[61] =16'd1563 ;
			a[62] =16'd34498;
			a[63] =16'd35617;
			temp_mult[576] = mult[0] ;
			temp_mult[577] = mult[1] ;
			temp_mult[578] = mult[2] ;
			temp_mult[579] = mult[3] ;
			temp_mult[580] = mult[4] ;
			temp_mult[581] = mult[5] ;
			temp_mult[582] = mult[6] ;
			temp_mult[583] = mult[7] ;
			temp_mult[584] = mult[8] ;
			temp_mult[585] = mult[9] ;
			temp_mult[586] = mult[10];
			temp_mult[587] = mult[11];
			temp_mult[588] = mult[12];
			temp_mult[589] = mult[13];
			temp_mult[590] = mult[14];
			temp_mult[591] = mult[15];
			temp_mult[592] = mult[16];
			temp_mult[593] = mult[17];
			temp_mult[594] = mult[18];
			temp_mult[595] = mult[19];
			temp_mult[596] = mult[20];
			temp_mult[597] = mult[21];
			temp_mult[598] = mult[22];
			temp_mult[599] = mult[23];
			temp_mult[600] = mult[24];
			temp_mult[601] = mult[25];
			temp_mult[602] = mult[26];
			temp_mult[603] = mult[27];
			temp_mult[604] = mult[28];
			temp_mult[605] = mult[29];
			temp_mult[606] = mult[30];
			temp_mult[607] = mult[31];
			temp_mult[608] = mult[32];
			temp_mult[609] = mult[33];
			temp_mult[610] = mult[34];
			temp_mult[611] = mult[35];
			temp_mult[612] = mult[36];
			temp_mult[613] = mult[37];
			temp_mult[614] = mult[38];
			temp_mult[615] = mult[39];
			temp_mult[616] = mult[40];
			temp_mult[617] = mult[41];
			temp_mult[618] = mult[42];
			temp_mult[619] = mult[43];
			temp_mult[620] = mult[44];
			temp_mult[621] = mult[45];
			temp_mult[622] = mult[46];
			temp_mult[623] = mult[47];
			temp_mult[624] = mult[48];
			temp_mult[625] = mult[49];
			temp_mult[626] = mult[50];
			temp_mult[627] = mult[51];
			temp_mult[628] = mult[52];
			temp_mult[629] = mult[53];
			temp_mult[630] = mult[54];
			temp_mult[631] = mult[55];
			temp_mult[632] = mult[56];
			temp_mult[633] = mult[57];
			temp_mult[634] = mult[58];
			temp_mult[635] = mult[59];
			temp_mult[636] = mult[60];
			temp_mult[637] = mult[61];
			temp_mult[638] = mult[62];
			temp_mult[639] = mult[63];
		end
		5'd11: begin
			b[0]  = d1_input_r[128];
			b[1]  = d1_input_r[129];
			b[2]  = d1_input_r[130];
			b[3]  = d1_input_r[131];
			b[4]  = d1_input_r[132];
			b[5]  = d1_input_r[133];
			b[6]  = d1_input_r[134];
			b[7]  = d1_input_r[135];
			b[8]  = d1_input_r[136];
			b[9]  = d1_input_r[137];
			b[10] = d1_input_r[138];
			b[11] = d1_input_r[139];
			b[12] = d1_input_r[140];
			b[13] = d1_input_r[141];
			b[14] = d1_input_r[142];
			b[15] = d1_input_r[143];
			b[16] = d1_input_r[144];
			b[17] = d1_input_r[145];
			b[18] = d1_input_r[146];
			b[19] = d1_input_r[147];
			b[20] = d1_input_r[148];
			b[21] = d1_input_r[149];
			b[22] = d1_input_r[150];
			b[23] = d1_input_r[151];
			b[24] = d1_input_r[152];
			b[25] = d1_input_r[153];
			b[26] = d1_input_r[154];
			b[27] = d1_input_r[155];
			b[28] = d1_input_r[156];
			b[29] = d1_input_r[157];
			b[30] = d1_input_r[158];
			b[31] = d1_input_r[159];
			b[32] = d1_input_r[160];
			b[33] = d1_input_r[161];
			b[34] = d1_input_r[162];
			b[35] = d1_input_r[163];
			b[36] = d1_input_r[164];
			b[37] = d1_input_r[165];
			b[38] = d1_input_r[166];
			b[39] = d1_input_r[167];
			b[40] = d1_input_r[168];
			b[41] = d1_input_r[169];
			b[42] = d1_input_r[170];
			b[43] = d1_input_r[171];
			b[44] = d1_input_r[172];
			b[45] = d1_input_r[173];
			b[46] = d1_input_r[174];
			b[47] = d1_input_r[175];
			b[48] = d1_input_r[176];
			b[49] = d1_input_r[177];
			b[50] = d1_input_r[178];
			b[51] = d1_input_r[179];
			b[52] = d1_input_r[180];
			b[53] = d1_input_r[181];
			b[54] = d1_input_r[182];
			b[55] = d1_input_r[183];
			b[56] = d1_input_r[184];
			b[57] = d1_input_r[185];
			b[58] = d1_input_r[186];
			b[59] = d1_input_r[187];
			b[60] = d1_input_r[188];
			b[61] = d1_input_r[189];
			b[62] = d1_input_r[190];
			b[63] = d1_input_r[191];
			a[0]  =16'd33841;
			a[1]  =16'd1287 ;
			a[2]  =16'd1636 ;
			a[3]  =16'd34680;
			a[4]  =16'd1541 ;
			a[5]  =16'd1766 ;
			a[6]  =16'd1920 ;
			a[7]  =16'd35818;
			a[8]  =16'd1451 ;
			a[9]  =16'd2417 ;
			a[10] =16'd34665;
			a[11] =16'd2462 ;
			a[12] =16'd33322;
			a[13] =16'd35852;
			a[14] =16'd33083;
			a[15] =16'd32940;
			a[16] =16'd1868 ;
			a[17] =16'd35512;
			a[18] =16'd33088;
			a[19] =16'd33373;
			a[20] =16'd32838;
			a[21] =16'd33159;
			a[22] =16'd225  ;
			a[23] =16'd1899 ;
			a[24] =16'd33463;
			a[25] =16'd264  ;
			a[26] =16'd33642;
			a[27] =16'd33501;
			a[28] =16'd1393 ;
			a[29] =16'd34539;
			a[30] =16'd32901;
			a[31] =16'd34254;
			a[32] =16'd33101;
			a[33] =16'd33289;
			a[34] =16'd34653;
			a[35] =16'd32795;
			a[36] =16'd35440;
			a[37] =16'd33852;
			a[38] =16'd756  ;
			a[39] =16'd35268;
			a[40] =16'd1808 ;
			a[41] =16'd33602;
			a[42] =16'd1456 ;
			a[43] =16'd32960;
			a[44] =16'd34305;
			a[45] =16'd955  ;
			a[46] =16'd32814;
			a[47] =16'd1790 ;
			a[48] =16'd404  ;
			a[49] =16'd33401;
			a[50] =16'd598  ;
			a[51] =16'd34933;
			a[52] =16'd34034;
			a[53] =16'd2652 ;
			a[54] =16'd1940 ;
			a[55] =16'd33622;
			a[56] =16'd34213;
			a[57] =16'd32877;
			a[58] =16'd34691;
			a[59] =16'd1503 ;
			a[60] =16'd1608 ;
			a[61] =16'd34270;
			a[62] =16'd508  ;
			a[63] =16'd35404;
			temp_mult[640] = mult[0] ;
			temp_mult[641] = mult[1] ;
			temp_mult[642] = mult[2] ;
			temp_mult[643] = mult[3] ;
			temp_mult[644] = mult[4] ;
			temp_mult[645] = mult[5] ;
			temp_mult[646] = mult[6] ;
			temp_mult[647] = mult[7] ;
			temp_mult[648] = mult[8] ;
			temp_mult[649] = mult[9] ;
			temp_mult[650] = mult[10];
			temp_mult[651] = mult[11];
			temp_mult[652] = mult[12];
			temp_mult[653] = mult[13];
			temp_mult[654] = mult[14];
			temp_mult[655] = mult[15];
			temp_mult[656] = mult[16];
			temp_mult[657] = mult[17];
			temp_mult[658] = mult[18];
			temp_mult[659] = mult[19];
			temp_mult[660] = mult[20];
			temp_mult[661] = mult[21];
			temp_mult[662] = mult[22];
			temp_mult[663] = mult[23];
			temp_mult[664] = mult[24];
			temp_mult[665] = mult[25];
			temp_mult[666] = mult[26];
			temp_mult[667] = mult[27];
			temp_mult[668] = mult[28];
			temp_mult[669] = mult[29];
			temp_mult[670] = mult[30];
			temp_mult[671] = mult[31];
			temp_mult[672] = mult[32];
			temp_mult[673] = mult[33];
			temp_mult[674] = mult[34];
			temp_mult[675] = mult[35];
			temp_mult[676] = mult[36];
			temp_mult[677] = mult[37];
			temp_mult[678] = mult[38];
			temp_mult[679] = mult[39];
			temp_mult[680] = mult[40];
			temp_mult[681] = mult[41];
			temp_mult[682] = mult[42];
			temp_mult[683] = mult[43];
			temp_mult[684] = mult[44];
			temp_mult[685] = mult[45];
			temp_mult[686] = mult[46];
			temp_mult[687] = mult[47];
			temp_mult[688] = mult[48];
			temp_mult[689] = mult[49];
			temp_mult[690] = mult[50];
			temp_mult[691] = mult[51];
			temp_mult[692] = mult[52];
			temp_mult[693] = mult[53];
			temp_mult[694] = mult[54];
			temp_mult[695] = mult[55];
			temp_mult[696] = mult[56];
			temp_mult[697] = mult[57];
			temp_mult[698] = mult[58];
			temp_mult[699] = mult[59];
			temp_mult[700] = mult[60];
			temp_mult[701] = mult[61];
			temp_mult[702] = mult[62];
			temp_mult[703] = mult[63];
		end
		5'd12: begin
			b[0]  = d1_input_r[192];
			b[1]  = d1_input_r[193];
			b[2]  = d1_input_r[194];
			b[3]  = d1_input_r[195];
			b[4]  = d1_input_r[196];
			b[5]  = d1_input_r[197];
			b[6]  = d1_input_r[198];
			b[7]  = d1_input_r[199];
			b[8]  = d1_input_r[200];
			b[9]  = d1_input_r[201];
			b[10] = d1_input_r[202];
			b[11] = d1_input_r[203];
			b[12] = d1_input_r[204];
			b[13] = d1_input_r[205];
			b[14] = d1_input_r[206];
			b[15] = d1_input_r[207];
			b[16] = d1_input_r[208];
			b[17] = d1_input_r[209];
			b[18] = d1_input_r[210];
			b[19] = d1_input_r[211];
			b[20] = d1_input_r[212];
			b[21] = d1_input_r[213];
			b[22] = d1_input_r[214];
			b[23] = d1_input_r[215];
			b[24] = d1_input_r[216];
			b[25] = d1_input_r[217];
			b[26] = d1_input_r[218];
			b[27] = d1_input_r[219];
			b[28] = d1_input_r[220];
			b[29] = d1_input_r[221];
			b[30] = d1_input_r[222];
			b[31] = d1_input_r[223];
			b[32] = d1_input_r[224];
			b[33] = d1_input_r[225];
			b[34] = d1_input_r[226];
			b[35] = d1_input_r[227];
			b[36] = d1_input_r[228];
			b[37] = d1_input_r[229];
			b[38] = d1_input_r[230];
			b[39] = d1_input_r[231];
			b[40] = d1_input_r[232];
			b[41] = d1_input_r[233];
			b[42] = d1_input_r[234];
			b[43] = d1_input_r[235];
			b[44] = d1_input_r[236];
			b[45] = d1_input_r[237];
			b[46] = d1_input_r[238];
			b[47] = d1_input_r[239];
			b[48] = d1_input_r[240];
			b[49] = d1_input_r[241];
			b[50] = d1_input_r[242];
			b[51] = d1_input_r[243];
			b[52] = d1_input_r[244];
			b[53] = d1_input_r[245];
			b[54] = d1_input_r[246];
			b[55] = d1_input_r[247];
			b[56] = d1_input_r[248];
			b[57] = d1_input_r[249];
			b[58] = d1_input_r[250];
			b[59] = d1_input_r[251];
			b[60] = d1_input_r[252];
			b[61] = d1_input_r[253];
			b[62] = d1_input_r[254];
			b[63] = d1_input_r[255];
			a[0]  =16'd34417;
			a[1]  =16'd973  ;
			a[2]  =16'd35455;
			a[3]  =16'd33200;
			a[4]  =16'd34772;
			a[5]  =16'd335  ;
			a[6]  =16'd33776;
			a[7]  =16'd1079 ;
			a[8]  =16'd34333;
			a[9]  =16'd33480;
			a[10] =16'd33876;
			a[11] =16'd110  ;
			a[12] =16'd35795;
			a[13] =16'd35338;
			a[14] =16'd34021;
			a[15] =16'd2448 ;
			a[16] =16'd2575 ;
			a[17] =16'd1248 ;
			a[18] =16'd1278 ;
			a[19] =16'd574  ;
			a[20] =16'd1197 ;
			a[21] =16'd2244 ;
			a[22] =16'd671  ;
			a[23] =16'd32774;
			a[24] =16'd883  ;
			a[25] =16'd914  ;
			a[26] =16'd35121;
			a[27] =16'd534  ;
			a[28] =16'd32856;
			a[29] =16'd33641;
			a[30] =16'd786  ;
			a[31] =16'd44   ;
			a[32] =16'd35437;
			a[33] =16'd1231 ;
			a[34] =16'd2247 ;
			a[35] =16'd1578 ;
			a[36] =16'd32935;
			a[37] =16'd33113;
			a[38] =16'd33153;
			a[39] =16'd1108 ;
			a[40] =16'd34843;
			a[41] =16'd625  ;
			a[42] =16'd2587 ;
			a[43] =16'd34189;
			a[44] =16'd2606 ;
			a[45] =16'd34205;
			a[46] =16'd33968;
			a[47] =16'd2741 ;
			a[48] =16'd1787 ;
			a[49] =16'd34089;
			a[50] =16'd33357;
			a[51] =16'd35082;
			a[52] =16'd413  ;
			a[53] =16'd34451;
			a[54] =16'd813  ;
			a[55] =16'd35048;
			a[56] =16'd34781;
			a[57] =16'd2325 ;
			a[58] =16'd32962;
			a[59] =16'd33548;
			a[60] =16'd728  ;
			a[61] =16'd1957 ;
			a[62] =16'd33473;
			a[63] =16'd35034;
			temp_mult[704] = mult[0] ;
			temp_mult[705] = mult[1] ;
			temp_mult[706] = mult[2] ;
			temp_mult[707] = mult[3] ;
			temp_mult[708] = mult[4] ;
			temp_mult[709] = mult[5] ;
			temp_mult[710] = mult[6] ;
			temp_mult[711] = mult[7] ;
			temp_mult[712] = mult[8] ;
			temp_mult[713] = mult[9] ;
			temp_mult[714] = mult[10];
			temp_mult[715] = mult[11];
			temp_mult[716] = mult[12];
			temp_mult[717] = mult[13];
			temp_mult[718] = mult[14];
			temp_mult[719] = mult[15];
			temp_mult[720] = mult[16];
			temp_mult[721] = mult[17];
			temp_mult[722] = mult[18];
			temp_mult[723] = mult[19];
			temp_mult[724] = mult[20];
			temp_mult[725] = mult[21];
			temp_mult[726] = mult[22];
			temp_mult[727] = mult[23];
			temp_mult[728] = mult[24];
			temp_mult[729] = mult[25];
			temp_mult[730] = mult[26];
			temp_mult[731] = mult[27];
			temp_mult[732] = mult[28];
			temp_mult[733] = mult[29];
			temp_mult[734] = mult[30];
			temp_mult[735] = mult[31];
			temp_mult[736] = mult[32];
			temp_mult[737] = mult[33];
			temp_mult[738] = mult[34];
			temp_mult[739] = mult[35];
			temp_mult[740] = mult[36];
			temp_mult[741] = mult[37];
			temp_mult[742] = mult[38];
			temp_mult[743] = mult[39];
			temp_mult[744] = mult[40];
			temp_mult[745] = mult[41];
			temp_mult[746] = mult[42];
			temp_mult[747] = mult[43];
			temp_mult[748] = mult[44];
			temp_mult[749] = mult[45];
			temp_mult[750] = mult[46];
			temp_mult[751] = mult[47];
			temp_mult[752] = mult[48];
			temp_mult[753] = mult[49];
			temp_mult[754] = mult[50];
			temp_mult[755] = mult[51];
			temp_mult[756] = mult[52];
			temp_mult[757] = mult[53];
			temp_mult[758] = mult[54];
			temp_mult[759] = mult[55];
			temp_mult[760] = mult[56];
			temp_mult[761] = mult[57];
			temp_mult[762] = mult[58];
			temp_mult[763] = mult[59];
			temp_mult[764] = mult[60];
			temp_mult[765] = mult[61];
			temp_mult[766] = mult[62];
			temp_mult[767] = mult[63];
		end
		5'd13: begin
			b[0]  =  d1_input_r[0];
			b[1]  =  d1_input_r[1];
			b[2]  =  d1_input_r[2];
			b[3]  =  d1_input_r[3];
			b[4]  =  d1_input_r[4];
			b[5]  =  d1_input_r[5];
			b[6]  =  d1_input_r[6];
			b[7]  =  d1_input_r[7];
			b[8]  =  d1_input_r[8];
			b[9]  =  d1_input_r[9];
			b[10] =  d1_input_r[10];
			b[11] =  d1_input_r[11];
			b[12] =  d1_input_r[12];
			b[13] =  d1_input_r[13];
			b[14] =  d1_input_r[14];
			b[15] =  d1_input_r[15];
			b[16] =  d1_input_r[16];
			b[17] =  d1_input_r[17];
			b[18] =  d1_input_r[18];
			b[19] =  d1_input_r[19];
			b[20] =  d1_input_r[20];
			b[21] =  d1_input_r[21];
			b[22] =  d1_input_r[22];
			b[23] =  d1_input_r[23];
			b[24] =  d1_input_r[24];
			b[25] =  d1_input_r[25];
			b[26] =  d1_input_r[26];
			b[27] =  d1_input_r[27];
			b[28] =  d1_input_r[28];
			b[29] =  d1_input_r[29];
			b[30] =  d1_input_r[30];
			b[31] =  d1_input_r[31];
			b[32] =  d1_input_r[32];
			b[33] =  d1_input_r[33];
			b[34] =  d1_input_r[34];
			b[35] =  d1_input_r[35];
			b[36] =  d1_input_r[36];
			b[37] =  d1_input_r[37];
			b[38] =  d1_input_r[38];
			b[39] =  d1_input_r[39];
			b[40] =  d1_input_r[40];
			b[41] =  d1_input_r[41];
			b[42] =  d1_input_r[42];
			b[43] =  d1_input_r[43];
			b[44] =  d1_input_r[44];
			b[45] =  d1_input_r[45];
			b[46] =  d1_input_r[46];
			b[47] =  d1_input_r[47];
			b[48] =  d1_input_r[48];
			b[49] =  d1_input_r[49];
			b[50] =  d1_input_r[50];
			b[51] =  d1_input_r[51];
			b[52] =  d1_input_r[52];
			b[53] =  d1_input_r[53];
			b[54] =  d1_input_r[54];
			b[55] =  d1_input_r[55];
			b[56] =  d1_input_r[56];
			b[57] =  d1_input_r[57];
			b[58] =  d1_input_r[58];
			b[59] =  d1_input_r[59];
			b[60] =  d1_input_r[60];
			b[61] =  d1_input_r[61];
			b[62] =  d1_input_r[62];
			b[63] =  d1_input_r[63];
			a[0]  =16'd34438;
			a[1]  =16'd341  ;
			a[2]  =16'd2510 ;
			a[3]  =16'd35385;
			a[4]  =16'd33538;
			a[5]  =16'd1219 ;
			a[6]  =16'd34335;
			a[7]  =16'd359  ;
			a[8]  =16'd33769;
			a[9]  =16'd785  ;
			a[10] =16'd795  ;
			a[11] =16'd34594;
			a[12] =16'd32802;
			a[13] =16'd218  ;
			a[14] =16'd35876;
			a[15] =16'd34609;
			a[16] =16'd33842;
			a[17] =16'd2030 ;
			a[18] =16'd1441 ;
			a[19] =16'd1348 ;
			a[20] =16'd2549 ;
			a[21] =16'd143  ;
			a[22] =16'd32903;
			a[23] =16'd893  ;
			a[24] =16'd33551;
			a[25] =16'd32940;
			a[26] =16'd33418;
			a[27] =16'd33002;
			a[28] =16'd1182 ;
			a[29] =16'd2320 ;
			a[30] =16'd33257;
			a[31] =16'd34917;
			a[32] =16'd34833;
			a[33] =16'd1530 ;
			a[34] =16'd33458;
			a[35] =16'd34845;
			a[36] =16'd34334;
			a[37] =16'd71   ;
			a[38] =16'd750  ;
			a[39] =16'd34882;
			a[40] =16'd315  ;
			a[41] =16'd34564;
			a[42] =16'd33520;
			a[43] =16'd34593;
			a[44] =16'd33381;
			a[45] =16'd1810 ;
			a[46] =16'd2352 ;
			a[47] =16'd2566 ;
			a[48] =16'd33629;
			a[49] =16'd420  ;
			a[50] =16'd2279 ;
			a[51] =16'd33448;
			a[52] =16'd34339;
			a[53] =16'd35377;
			a[54] =16'd1390 ;
			a[55] =16'd1097 ;
			a[56] =16'd1419 ;
			a[57] =16'd35001;
			a[58] =16'd3022 ;
			a[59] =16'd35292;
			a[60] =16'd35208;
			a[61] =16'd34584;
			a[62] =16'd2189 ;
			a[63] =16'd33479;
			temp_mult[768] = mult[0] ;
			temp_mult[769] = mult[1] ;
			temp_mult[770] = mult[2] ;
			temp_mult[771] = mult[3] ;
			temp_mult[772] = mult[4] ;
			temp_mult[773] = mult[5] ;
			temp_mult[774] = mult[6] ;
			temp_mult[775] = mult[7] ;
			temp_mult[776] = mult[8] ;
			temp_mult[777] = mult[9] ;
			temp_mult[778] = mult[10];
			temp_mult[779] = mult[11];
			temp_mult[780] = mult[12];
			temp_mult[781] = mult[13];
			temp_mult[782] = mult[14];
			temp_mult[783] = mult[15];
			temp_mult[784] = mult[16];
			temp_mult[785] = mult[17];
			temp_mult[786] = mult[18];
			temp_mult[787] = mult[19];
			temp_mult[788] = mult[20];
			temp_mult[789] = mult[21];
			temp_mult[790] = mult[22];
			temp_mult[791] = mult[23];
			temp_mult[792] = mult[24];
			temp_mult[793] = mult[25];
			temp_mult[794] = mult[26];
			temp_mult[795] = mult[27];
			temp_mult[796] = mult[28];
			temp_mult[797] = mult[29];
			temp_mult[798] = mult[30];
			temp_mult[799] = mult[31];
			temp_mult[800] = mult[32];
			temp_mult[801] = mult[33];
			temp_mult[802] = mult[34];
			temp_mult[803] = mult[35];
			temp_mult[804] = mult[36];
			temp_mult[805] = mult[37];
			temp_mult[806] = mult[38];
			temp_mult[807] = mult[39];
			temp_mult[808] = mult[40];
			temp_mult[809] = mult[41];
			temp_mult[810] = mult[42];
			temp_mult[811] = mult[43];
			temp_mult[812] = mult[44];
			temp_mult[813] = mult[45];
			temp_mult[814] = mult[46];
			temp_mult[815] = mult[47];
			temp_mult[816] = mult[48];
			temp_mult[817] = mult[49];
			temp_mult[818] = mult[50];
			temp_mult[819] = mult[51];
			temp_mult[820] = mult[52];
			temp_mult[821] = mult[53];
			temp_mult[822] = mult[54];
			temp_mult[823] = mult[55];
			temp_mult[824] = mult[56];
			temp_mult[825] = mult[57];
			temp_mult[826] = mult[58];
			temp_mult[827] = mult[59];
			temp_mult[828] = mult[60];
			temp_mult[829] = mult[61];
			temp_mult[830] = mult[62];
			temp_mult[831] = mult[63];
		end
		5'd14: begin
			b[0]  = d1_input_r[64];
			b[1]  = d1_input_r[65];
			b[2]  = d1_input_r[66];
			b[3]  = d1_input_r[67];
			b[4]  = d1_input_r[68];
			b[5]  = d1_input_r[69];
			b[6]  = d1_input_r[70];
			b[7]  = d1_input_r[71];
			b[8]  = d1_input_r[72];
			b[9]  = d1_input_r[73];
			b[10] = d1_input_r[74];
			b[11] = d1_input_r[75];
			b[12] = d1_input_r[76];
			b[13] = d1_input_r[77];
			b[14] = d1_input_r[78];
			b[15] = d1_input_r[79];
			b[16] = d1_input_r[80];
			b[17] = d1_input_r[81];
			b[18] = d1_input_r[82];
			b[19] = d1_input_r[83];
			b[20] = d1_input_r[84];
			b[21] = d1_input_r[85];
			b[22] = d1_input_r[86];
			b[23] = d1_input_r[87];
			b[24] = d1_input_r[88];
			b[25] = d1_input_r[89];
			b[26] = d1_input_r[90];
			b[27] = d1_input_r[91];
			b[28] = d1_input_r[92];
			b[29] = d1_input_r[93];
			b[30] = d1_input_r[94];
			b[31] = d1_input_r[95];
			b[32] = d1_input_r[96];
			b[33] = d1_input_r[97];
			b[34] = d1_input_r[98];
			b[35] = d1_input_r[99];
			b[36] = d1_input_r[100];
			b[37] = d1_input_r[101];
			b[38] = d1_input_r[102];
			b[39] = d1_input_r[103];
			b[40] = d1_input_r[104];
			b[41] = d1_input_r[105];
			b[42] = d1_input_r[106];
			b[43] = d1_input_r[107];
			b[44] = d1_input_r[108];
			b[45] = d1_input_r[109];
			b[46] = d1_input_r[110];
			b[47] = d1_input_r[111];
			b[48] = d1_input_r[112];
			b[49] = d1_input_r[113];
			b[50] = d1_input_r[114];
			b[51] = d1_input_r[115];
			b[52] = d1_input_r[116];
			b[53] = d1_input_r[117];
			b[54] = d1_input_r[118];
			b[55] = d1_input_r[119];
			b[56] = d1_input_r[120];
			b[57] = d1_input_r[121];
			b[58] = d1_input_r[122];
			b[59] = d1_input_r[123];
			b[60] = d1_input_r[124];
			b[61] = d1_input_r[125];
			b[62] = d1_input_r[126];
			b[63] = d1_input_r[127];
			a[0]  =16'd35315;
			a[1]  =16'd836  ;
			a[2]  =16'd2041 ;
			a[3]  =16'd35457;
			a[4]  =16'd1651 ;
			a[5]  =16'd828  ;
			a[6]  =16'd872  ;
			a[7]  =16'd539  ;
			a[8]  =16'd1319 ;
			a[9]  =16'd34557;
			a[10] =16'd33301;
			a[11] =16'd579  ;
			a[12] =16'd33173;
			a[13] =16'd334  ;
			a[14] =16'd2210 ;
			a[15] =16'd2884 ;
			a[16] =16'd1616 ;
			a[17] =16'd33196;
			a[18] =16'd873  ;
			a[19] =16'd33970;
			a[20] =16'd1410 ;
			a[21] =16'd34550;
			a[22] =16'd34430;
			a[23] =16'd33926;
			a[24] =16'd35229;
			a[25] =16'd2849 ;
			a[26] =16'd801  ;
			a[27] =16'd34141;
			a[28] =16'd33958;
			a[29] =16'd2924 ;
			a[30] =16'd1920 ;
			a[31] =16'd35771;
			a[32] =16'd1843 ;
			a[33] =16'd513  ;
			a[34] =16'd33657;
			a[35] =16'd35732;
			a[36] =16'd2142 ;
			a[37] =16'd2260 ;
			a[38] =16'd2037 ;
			a[39] =16'd33969;
			a[40] =16'd35041;
			a[41] =16'd2275 ;
			a[42] =16'd354  ;
			a[43] =16'd34734;
			a[44] =16'd122  ;
			a[45] =16'd1517 ;
			a[46] =16'd1969 ;
			a[47] =16'd32775;
			a[48] =16'd33170;
			a[49] =16'd34598;
			a[50] =16'd34679;
			a[51] =16'd33162;
			a[52] =16'd554  ;
			a[53] =16'd34034;
			a[54] =16'd33987;
			a[55] =16'd1250 ;
			a[56] =16'd32908;
			a[57] =16'd33551;
			a[58] =16'd1151 ;
			a[59] =16'd35741;
			a[60] =16'd1221 ;
			a[61] =16'd34138;
			a[62] =16'd1526 ;
			a[63] =16'd1135 ;
			temp_mult[832] = mult[0] ;
			temp_mult[833] = mult[1] ;
			temp_mult[834] = mult[2] ;
			temp_mult[835] = mult[3] ;
			temp_mult[836] = mult[4] ;
			temp_mult[837] = mult[5] ;
			temp_mult[838] = mult[6] ;
			temp_mult[839] = mult[7] ;
			temp_mult[840] = mult[8] ;
			temp_mult[841] = mult[9] ;
			temp_mult[842] = mult[10];
			temp_mult[843] = mult[11];
			temp_mult[844] = mult[12];
			temp_mult[845] = mult[13];
			temp_mult[846] = mult[14];
			temp_mult[847] = mult[15];
			temp_mult[848] = mult[16];
			temp_mult[849] = mult[17];
			temp_mult[850] = mult[18];
			temp_mult[851] = mult[19];
			temp_mult[852] = mult[20];
			temp_mult[853] = mult[21];
			temp_mult[854] = mult[22];
			temp_mult[855] = mult[23];
			temp_mult[856] = mult[24];
			temp_mult[857] = mult[25];
			temp_mult[858] = mult[26];
			temp_mult[859] = mult[27];
			temp_mult[860] = mult[28];
			temp_mult[861] = mult[29];
			temp_mult[862] = mult[30];
			temp_mult[863] = mult[31];
			temp_mult[864] = mult[32];
			temp_mult[865] = mult[33];
			temp_mult[866] = mult[34];
			temp_mult[867] = mult[35];
			temp_mult[868] = mult[36];
			temp_mult[869] = mult[37];
			temp_mult[870] = mult[38];
			temp_mult[871] = mult[39];
			temp_mult[872] = mult[40];
			temp_mult[873] = mult[41];
			temp_mult[874] = mult[42];
			temp_mult[875] = mult[43];
			temp_mult[876] = mult[44];
			temp_mult[877] = mult[45];
			temp_mult[878] = mult[46];
			temp_mult[879] = mult[47];
			temp_mult[880] = mult[48];
			temp_mult[881] = mult[49];
			temp_mult[882] = mult[50];
			temp_mult[883] = mult[51];
			temp_mult[884] = mult[52];
			temp_mult[885] = mult[53];
			temp_mult[886] = mult[54];
			temp_mult[887] = mult[55];
			temp_mult[888] = mult[56];
			temp_mult[889] = mult[57];
			temp_mult[890] = mult[58];
			temp_mult[891] = mult[59];
			temp_mult[892] = mult[60];
			temp_mult[893] = mult[61];
			temp_mult[894] = mult[62];
			temp_mult[895] = mult[63];
		end
		5'd15: begin
			b[0]  = d1_input_r[128];
			b[1]  = d1_input_r[129];
			b[2]  = d1_input_r[130];
			b[3]  = d1_input_r[131];
			b[4]  = d1_input_r[132];
			b[5]  = d1_input_r[133];
			b[6]  = d1_input_r[134];
			b[7]  = d1_input_r[135];
			b[8]  = d1_input_r[136];
			b[9]  = d1_input_r[137];
			b[10] = d1_input_r[138];
			b[11] = d1_input_r[139];
			b[12] = d1_input_r[140];
			b[13] = d1_input_r[141];
			b[14] = d1_input_r[142];
			b[15] = d1_input_r[143];
			b[16] = d1_input_r[144];
			b[17] = d1_input_r[145];
			b[18] = d1_input_r[146];
			b[19] = d1_input_r[147];
			b[20] = d1_input_r[148];
			b[21] = d1_input_r[149];
			b[22] = d1_input_r[150];
			b[23] = d1_input_r[151];
			b[24] = d1_input_r[152];
			b[25] = d1_input_r[153];
			b[26] = d1_input_r[154];
			b[27] = d1_input_r[155];
			b[28] = d1_input_r[156];
			b[29] = d1_input_r[157];
			b[30] = d1_input_r[158];
			b[31] = d1_input_r[159];
			b[32] = d1_input_r[160];
			b[33] = d1_input_r[161];
			b[34] = d1_input_r[162];
			b[35] = d1_input_r[163];
			b[36] = d1_input_r[164];
			b[37] = d1_input_r[165];
			b[38] = d1_input_r[166];
			b[39] = d1_input_r[167];
			b[40] = d1_input_r[168];
			b[41] = d1_input_r[169];
			b[42] = d1_input_r[170];
			b[43] = d1_input_r[171];
			b[44] = d1_input_r[172];
			b[45] = d1_input_r[173];
			b[46] = d1_input_r[174];
			b[47] = d1_input_r[175];
			b[48] = d1_input_r[176];
			b[49] = d1_input_r[177];
			b[50] = d1_input_r[178];
			b[51] = d1_input_r[179];
			b[52] = d1_input_r[180];
			b[53] = d1_input_r[181];
			b[54] = d1_input_r[182];
			b[55] = d1_input_r[183];
			b[56] = d1_input_r[184];
			b[57] = d1_input_r[185];
			b[58] = d1_input_r[186];
			b[59] = d1_input_r[187];
			b[60] = d1_input_r[188];
			b[61] = d1_input_r[189];
			b[62] = d1_input_r[190];
			b[63] = d1_input_r[191];
			a[0]  =16'd35909;
			a[1]  =16'd1661 ;
			a[2]  =16'd33812;
			a[3]  =16'd34957;
			a[4]  =16'd2074 ;
			a[5]  =16'd1265 ;
			a[6]  =16'd1475 ;
			a[7]  =16'd1647 ;
			a[8]  =16'd447  ;
			a[9]  =16'd33853;
			a[10] =16'd2479 ;
			a[11] =16'd486  ;
			a[12] =16'd33967;
			a[13] =16'd33295;
			a[14] =16'd34128;
			a[15] =16'd994  ;
			a[16] =16'd2530 ;
			a[17] =16'd33961;
			a[18] =16'd34945;
			a[19] =16'd34327;
			a[20] =16'd2964 ;
			a[21] =16'd1666 ;
			a[22] =16'd1429 ;
			a[23] =16'd33167;
			a[24] =16'd34985;
			a[25] =16'd2347 ;
			a[26] =16'd33469;
			a[27] =16'd32852;
			a[28] =16'd222  ;
			a[29] =16'd2049 ;
			a[30] =16'd1790 ;
			a[31] =16'd680  ;
			a[32] =16'd34420;
			a[33] =16'd2229 ;
			a[34] =16'd679  ;
			a[35] =16'd1516 ;
			a[36] =16'd1727 ;
			a[37] =16'd2135 ;
			a[38] =16'd34397;
			a[39] =16'd33511;
			a[40] =16'd1000 ;
			a[41] =16'd33422;
			a[42] =16'd705  ;
			a[43] =16'd1811 ;
			a[44] =16'd33699;
			a[45] =16'd397  ;
			a[46] =16'd33596;
			a[47] =16'd433  ;
			a[48] =16'd33237;
			a[49] =16'd33933;
			a[50] =16'd34933;
			a[51] =16'd34687;
			a[52] =16'd2713 ;
			a[53] =16'd1122 ;
			a[54] =16'd33737;
			a[55] =16'd33743;
			a[56] =16'd793  ;
			a[57] =16'd2496 ;
			a[58] =16'd33328;
			a[59] =16'd803  ;
			a[60] =16'd33001;
			a[61] =16'd2735 ;
			a[62] =16'd1950 ;
			a[63] =16'd535  ;
			temp_mult[896] = mult[0] ;
			temp_mult[897] = mult[1] ;
			temp_mult[898] = mult[2] ;
			temp_mult[899] = mult[3] ;
			temp_mult[900] = mult[4] ;
			temp_mult[901] = mult[5] ;
			temp_mult[902] = mult[6] ;
			temp_mult[903] = mult[7] ;
			temp_mult[904] = mult[8] ;
			temp_mult[905] = mult[9] ;
			temp_mult[906] = mult[10];
			temp_mult[907] = mult[11];
			temp_mult[908] = mult[12];
			temp_mult[909] = mult[13];
			temp_mult[910] = mult[14];
			temp_mult[911] = mult[15];
			temp_mult[912] = mult[16];
			temp_mult[913] = mult[17];
			temp_mult[914] = mult[18];
			temp_mult[915] = mult[19];
			temp_mult[916] = mult[20];
			temp_mult[917] = mult[21];
			temp_mult[918] = mult[22];
			temp_mult[919] = mult[23];
			temp_mult[920] = mult[24];
			temp_mult[921] = mult[25];
			temp_mult[922] = mult[26];
			temp_mult[923] = mult[27];
			temp_mult[924] = mult[28];
			temp_mult[925] = mult[29];
			temp_mult[926] = mult[30];
			temp_mult[927] = mult[31];
			temp_mult[928] = mult[32];
			temp_mult[929] = mult[33];
			temp_mult[930] = mult[34];
			temp_mult[931] = mult[35];
			temp_mult[932] = mult[36];
			temp_mult[933] = mult[37];
			temp_mult[934] = mult[38];
			temp_mult[935] = mult[39];
			temp_mult[936] = mult[40];
			temp_mult[937] = mult[41];
			temp_mult[938] = mult[42];
			temp_mult[939] = mult[43];
			temp_mult[940] = mult[44];
			temp_mult[941] = mult[45];
			temp_mult[942] = mult[46];
			temp_mult[943] = mult[47];
			temp_mult[944] = mult[48];
			temp_mult[945] = mult[49];
			temp_mult[946] = mult[50];
			temp_mult[947] = mult[51];
			temp_mult[948] = mult[52];
			temp_mult[949] = mult[53];
			temp_mult[950] = mult[54];
			temp_mult[951] = mult[55];
			temp_mult[952] = mult[56];
			temp_mult[953] = mult[57];
			temp_mult[954] = mult[58];
			temp_mult[955] = mult[59];
			temp_mult[956] = mult[60];
			temp_mult[957] = mult[61];
			temp_mult[958] = mult[62];
			temp_mult[959] = mult[63];
		end
		5'd16: begin
			b[0]  = d1_input_r[192];
			b[1]  = d1_input_r[193];
			b[2]  = d1_input_r[194];
			b[3]  = d1_input_r[195];
			b[4]  = d1_input_r[196];
			b[5]  = d1_input_r[197];
			b[6]  = d1_input_r[198];
			b[7]  = d1_input_r[199];
			b[8]  = d1_input_r[200];
			b[9]  = d1_input_r[201];
			b[10] = d1_input_r[202];
			b[11] = d1_input_r[203];
			b[12] = d1_input_r[204];
			b[13] = d1_input_r[205];
			b[14] = d1_input_r[206];
			b[15] = d1_input_r[207];
			b[16] = d1_input_r[208];
			b[17] = d1_input_r[209];
			b[18] = d1_input_r[210];
			b[19] = d1_input_r[211];
			b[20] = d1_input_r[212];
			b[21] = d1_input_r[213];
			b[22] = d1_input_r[214];
			b[23] = d1_input_r[215];
			b[24] = d1_input_r[216];
			b[25] = d1_input_r[217];
			b[26] = d1_input_r[218];
			b[27] = d1_input_r[219];
			b[28] = d1_input_r[220];
			b[29] = d1_input_r[221];
			b[30] = d1_input_r[222];
			b[31] = d1_input_r[223];
			b[32] = d1_input_r[224];
			b[33] = d1_input_r[225];
			b[34] = d1_input_r[226];
			b[35] = d1_input_r[227];
			b[36] = d1_input_r[228];
			b[37] = d1_input_r[229];
			b[38] = d1_input_r[230];
			b[39] = d1_input_r[231];
			b[40] = d1_input_r[232];
			b[41] = d1_input_r[233];
			b[42] = d1_input_r[234];
			b[43] = d1_input_r[235];
			b[44] = d1_input_r[236];
			b[45] = d1_input_r[237];
			b[46] = d1_input_r[238];
			b[47] = d1_input_r[239];
			b[48] = d1_input_r[240];
			b[49] = d1_input_r[241];
			b[50] = d1_input_r[242];
			b[51] = d1_input_r[243];
			b[52] = d1_input_r[244];
			b[53] = d1_input_r[245];
			b[54] = d1_input_r[246];
			b[55] = d1_input_r[247];
			b[56] = d1_input_r[248];
			b[57] = d1_input_r[249];
			b[58] = d1_input_r[250];
			b[59] = d1_input_r[251];
			b[60] = d1_input_r[252];
			b[61] = d1_input_r[253];
			b[62] = d1_input_r[254];
			b[63] = d1_input_r[255];
			a[0]  =16'd35031;
			a[1]  =16'd1216 ;
			a[2]  =16'd34730;
			a[3]  =16'd32871;
			a[4]  =16'd802  ;
			a[5]  =16'd662  ;
			a[6]  =16'd33743;
			a[7]  =16'd516  ;
			a[8]  =16'd35665;
			a[9]  =16'd774  ;
			a[10] =16'd939  ;
			a[11] =16'd32816;
			a[12] =16'd34150;
			a[13] =16'd35420;
			a[14] =16'd1456 ;
			a[15] =16'd501  ;
			a[16] =16'd1190 ;
			a[17] =16'd34887;
			a[18] =16'd32966;
			a[19] =16'd34150;
			a[20] =16'd3008 ;
			a[21] =16'd34244;
			a[22] =16'd33623;
			a[23] =16'd1685 ;
			a[24] =16'd33213;
			a[25] =16'd2179 ;
			a[26] =16'd34125;
			a[27] =16'd1115 ;
			a[28] =16'd33935;
			a[29] =16'd2460 ;
			a[30] =16'd33038;
			a[31] =16'd33541;
			a[32] =16'd33742;
			a[33] =16'd1472 ;
			a[34] =16'd33436;
			a[35] =16'd1044 ;
			a[36] =16'd705  ;
			a[37] =16'd33431;
			a[38] =16'd34594;
			a[39] =16'd33268;
			a[40] =16'd34076;
			a[41] =16'd1060 ;
			a[42] =16'd32906;
			a[43] =16'd34681;
			a[44] =16'd33523;
			a[45] =16'd34134;
			a[46] =16'd1900 ;
			a[47] =16'd2208 ;
			a[48] =16'd1292 ;
			a[49] =16'd1152 ;
			a[50] =16'd35077;
			a[51] =16'd33308;
			a[52] =16'd34095;
			a[53] =16'd2222 ;
			a[54] =16'd34935;
			a[55] =16'd34745;
			a[56] =16'd34674;
			a[57] =16'd2328 ;
			a[58] =16'd34186;
			a[59] =16'd34893;
			a[60] =16'd35358;
			a[61] =16'd33389;
			a[62] =16'd291  ;
			a[63] =16'd35035;
			temp_mult[960] = mult[0] ;
			temp_mult[961] = mult[1] ;
			temp_mult[962] = mult[2] ;
			temp_mult[963] = mult[3] ;
			temp_mult[964] = mult[4] ;
			temp_mult[965] = mult[5] ;
			temp_mult[966] = mult[6] ;
			temp_mult[967] = mult[7] ;
			temp_mult[968] = mult[8] ;
			temp_mult[969] = mult[9] ;
			temp_mult[970] = mult[10];
			temp_mult[971] = mult[11];
			temp_mult[972] = mult[12];
			temp_mult[973] = mult[13];
			temp_mult[974] = mult[14];
			temp_mult[975] = mult[15];
			temp_mult[976] = mult[16];
			temp_mult[977] = mult[17];
			temp_mult[978] = mult[18];
			temp_mult[979] = mult[19];
			temp_mult[980] = mult[20];
			temp_mult[981] = mult[21];
			temp_mult[982] = mult[22];
			temp_mult[983] = mult[23];
			temp_mult[984] = mult[24];
			temp_mult[985] = mult[25];
			temp_mult[986] = mult[26];
			temp_mult[987] = mult[27];
			temp_mult[988] = mult[28];
			temp_mult[989] = mult[29];
			temp_mult[990] = mult[30];
			temp_mult[991] = mult[31];
			temp_mult[992] = mult[32];
			temp_mult[993] = mult[33];
			temp_mult[994] = mult[34];
			temp_mult[995] = mult[35];
			temp_mult[996] = mult[36];
			temp_mult[997] = mult[37];
			temp_mult[998] = mult[38];
			temp_mult[999] = mult[39];
			temp_mult[1000] = mult[40];
			temp_mult[1001] = mult[41];
			temp_mult[1002] = mult[42];
			temp_mult[1003] = mult[43];
			temp_mult[1004] = mult[44];
			temp_mult[1005] = mult[45];
			temp_mult[1006] = mult[46];
			temp_mult[1007] = mult[47];
			temp_mult[1008] = mult[48];
			temp_mult[1009] = mult[49];
			temp_mult[1010] = mult[50];
			temp_mult[1011] = mult[51];
			temp_mult[1012] = mult[52];
			temp_mult[1013] = mult[53];
			temp_mult[1014] = mult[54];
			temp_mult[1015] = mult[55];
			temp_mult[1016] = mult[56];
			temp_mult[1017] = mult[57];
			temp_mult[1018] = mult[58];
			temp_mult[1019] = mult[59];
			temp_mult[1020] = mult[60];
			temp_mult[1021] = mult[61];
			temp_mult[1022] = mult[62];
			temp_mult[1023] = mult[63];
		end
		default: begin
		
		end
	endcase
end

always @(*) begin
	if(!rst_n) begin
		temp_add[0] = 16'd0;
		temp_add[1] = 16'd0;
		temp_add[2] = 16'd0;
		temp_add[3] = 16'd0;
	end
	else begin
		for(i = 0; i < 256; i = i+1) begin
			temp_add[0] = temp_add[0] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
		for(i = 256; i < 512; i = i+1) begin
			temp_add[1] = temp_add[1] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
		for(i = 512; i < 768; i = i+1) begin
			temp_add[2] = temp_add[2] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
		for(i = 768; i < 1024; i = i+1) begin
			temp_add[3] = temp_add[3] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
	end
end

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		d1_output <= 64'd0;
		counter <= 5'd0;
	end
	else begin
		d1_output[15:0] <= temp_add[0] + bias[0];
		d1_output[31:16] <= temp_add[1] + bias[1];
		d1_output[47:32] <= temp_add[2] + bias[2];
		d1_output[63:48] <= temp_add[3] + bias[3];
		counter <= counter + 5'd1;
	end
end

endmodule