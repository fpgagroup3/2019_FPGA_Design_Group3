module	dense1(
	input clk,
	input rst_n,
	input [256*16-1:0] d1_input,
	output reg [4*16-1:0] d1_output
);


reg [15:0] d1_input_r [0:255];

wire [31:0] temp_mult [0:1023];
reg [15:0] temp_add [0:3];

wire [15:0] bias [0:3];

integer i, j;

assign bias[0] = 16'd346;
assign bias[1] = 16'd344; 
assign bias[2] = 16'd33106; 
assign bias[3] = 16'd33106;
assign temp_mult[0] = 16'd33087 * d1_input_r[0];
assign temp_mult[1] = 16'd198 * d1_input_r[1];
assign temp_mult[2] = 16'd34748 * d1_input_r[2];
assign temp_mult[3] = 16'd2210 * d1_input_r[3];
assign temp_mult[4] = 16'd1852 * d1_input_r[4];
assign temp_mult[5] = 16'd1435 * d1_input_r[5];
assign temp_mult[6] = 16'd157 * d1_input_r[6];
assign temp_mult[7] = 16'd1119 * d1_input_r[7];
assign temp_mult[8] = 16'd1120 * d1_input_r[8];
assign temp_mult[9] = 16'd986 * d1_input_r[9];
assign temp_mult[10] = 16'd1497 * d1_input_r[10];
assign temp_mult[11] = 16'd993 * d1_input_r[11];
assign temp_mult[12] = 16'd35132 * d1_input_r[12];
assign temp_mult[13] = 16'd2385 * d1_input_r[13];
assign temp_mult[14] = 16'd2952 * d1_input_r[14];
assign temp_mult[15] = 16'd35274 * d1_input_r[15];
assign temp_mult[16] = 16'd33781 * d1_input_r[16];
assign temp_mult[17] = 16'd1008 * d1_input_r[17];
assign temp_mult[18] = 16'd560 * d1_input_r[18];
assign temp_mult[19] = 16'd1522 * d1_input_r[19];
assign temp_mult[20] = 16'd33187 * d1_input_r[20];
assign temp_mult[21] = 16'd490 * d1_input_r[21];
assign temp_mult[22] = 16'd581 * d1_input_r[22];
assign temp_mult[23] = 16'd33711 * d1_input_r[23];
assign temp_mult[24] = 16'd32952 * d1_input_r[24];
assign temp_mult[25] = 16'd1612 * d1_input_r[25];
assign temp_mult[26] = 16'd948 * d1_input_r[26];
assign temp_mult[27] = 16'd94 * d1_input_r[27];
assign temp_mult[28] = 16'd32906 * d1_input_r[28];
assign temp_mult[29] = 16'd34931 * d1_input_r[29];
assign temp_mult[30] = 16'd33268 * d1_input_r[30];
assign temp_mult[31] = 16'd33834 * d1_input_r[31];
assign temp_mult[32] = 16'd138 * d1_input_r[32];
assign temp_mult[33] = 16'd33917 * d1_input_r[33];
assign temp_mult[34] = 16'd1104 * d1_input_r[34];
assign temp_mult[35] = 16'd34255 * d1_input_r[35];
assign temp_mult[36] = 16'd34349 * d1_input_r[36];
assign temp_mult[37] = 16'd33242 * d1_input_r[37];
assign temp_mult[38] = 16'd33852 * d1_input_r[38];
assign temp_mult[39] = 16'd717 * d1_input_r[39];
assign temp_mult[40] = 16'd1312 * d1_input_r[40];
assign temp_mult[41] = 16'd35246 * d1_input_r[41];
assign temp_mult[42] = 16'd2851 * d1_input_r[42];
assign temp_mult[43] = 16'd36 * d1_input_r[43];
assign temp_mult[44] = 16'd35195 * d1_input_r[44];
assign temp_mult[45] = 16'd35256 * d1_input_r[45];
assign temp_mult[46] = 16'd35134 * d1_input_r[46];
assign temp_mult[47] = 16'd1111 * d1_input_r[47];
assign temp_mult[48] = 16'd816 * d1_input_r[48];
assign temp_mult[49] = 16'd1649 * d1_input_r[49];
assign temp_mult[50] = 16'd33560 * d1_input_r[50];
assign temp_mult[51] = 16'd33982 * d1_input_r[51];
assign temp_mult[52] = 16'd1348 * d1_input_r[52];
assign temp_mult[53] = 16'd1352 * d1_input_r[53];
assign temp_mult[54] = 16'd870 * d1_input_r[54];
assign temp_mult[55] = 16'd1299 * d1_input_r[55];
assign temp_mult[56] = 16'd1142 * d1_input_r[56];
assign temp_mult[57] = 16'd33779 * d1_input_r[57];
assign temp_mult[58] = 16'd34197 * d1_input_r[58];
assign temp_mult[59] = 16'd174 * d1_input_r[59];
assign temp_mult[60] = 16'd2467 * d1_input_r[60];
assign temp_mult[61] = 16'd787 * d1_input_r[61];
assign temp_mult[62] = 16'd309 * d1_input_r[62];
assign temp_mult[63] = 16'd33043 * d1_input_r[63];
assign temp_mult[64] = 16'd33899 * d1_input_r[64];
assign temp_mult[65] = 16'd32983 * d1_input_r[65];
assign temp_mult[66] = 16'd2133 * d1_input_r[66];
assign temp_mult[67] = 16'd1803 * d1_input_r[67];
assign temp_mult[68] = 16'd1557 * d1_input_r[68];
assign temp_mult[69] = 16'd169 * d1_input_r[69];
assign temp_mult[70] = 16'd1054 * d1_input_r[70];
assign temp_mult[71] = 16'd1449 * d1_input_r[71];
assign temp_mult[72] = 16'd32910 * d1_input_r[72];
assign temp_mult[73] = 16'd34527 * d1_input_r[73];
assign temp_mult[74] = 16'd1212 * d1_input_r[74];
assign temp_mult[75] = 16'd1618 * d1_input_r[75];
assign temp_mult[76] = 16'd1457 * d1_input_r[76];
assign temp_mult[77] = 16'd563 * d1_input_r[77];
assign temp_mult[78] = 16'd33332 * d1_input_r[78];
assign temp_mult[79] = 16'd32956 * d1_input_r[79];
assign temp_mult[80] = 16'd1281 * d1_input_r[80];
assign temp_mult[81] = 16'd33648 * d1_input_r[81];
assign temp_mult[82] = 16'd1407 * d1_input_r[82];
assign temp_mult[83] = 16'd34453 * d1_input_r[83];
assign temp_mult[84] = 16'd35037 * d1_input_r[84];
assign temp_mult[85] = 16'd900 * d1_input_r[85];
assign temp_mult[86] = 16'd120 * d1_input_r[86];
assign temp_mult[87] = 16'd35796 * d1_input_r[87];
assign temp_mult[88] = 16'd34609 * d1_input_r[88];
assign temp_mult[89] = 16'd35377 * d1_input_r[89];
assign temp_mult[90] = 16'd1416 * d1_input_r[90];
assign temp_mult[91] = 16'd34359 * d1_input_r[91];
assign temp_mult[92] = 16'd2394 * d1_input_r[92];
assign temp_mult[93] = 16'd698 * d1_input_r[93];
assign temp_mult[94] = 16'd32824 * d1_input_r[94];
assign temp_mult[95] = 16'd33476 * d1_input_r[95];
assign temp_mult[96] = 16'd2785 * d1_input_r[96];
assign temp_mult[97] = 16'd33356 * d1_input_r[97];
assign temp_mult[98] = 16'd2651 * d1_input_r[98];
assign temp_mult[99] = 16'd33599 * d1_input_r[99];
assign temp_mult[100] = 16'd33773 * d1_input_r[100];
assign temp_mult[101] = 16'd726 * d1_input_r[101];
assign temp_mult[102] = 16'd1019 * d1_input_r[102];
assign temp_mult[103] = 16'd83 * d1_input_r[103];
assign temp_mult[104] = 16'd34379 * d1_input_r[104];
assign temp_mult[105] = 16'd34386 * d1_input_r[105];
assign temp_mult[106] = 16'd34448 * d1_input_r[106];
assign temp_mult[107] = 16'd33480 * d1_input_r[107];
assign temp_mult[108] = 16'd881 * d1_input_r[108];
assign temp_mult[109] = 16'd34240 * d1_input_r[109];
assign temp_mult[110] = 16'd1850 * d1_input_r[110];
assign temp_mult[111] = 16'd33793 * d1_input_r[111];
assign temp_mult[112] = 16'd33106 * d1_input_r[112];
assign temp_mult[113] = 16'd2276 * d1_input_r[113];
assign temp_mult[114] = 16'd33897 * d1_input_r[114];
assign temp_mult[115] = 16'd411 * d1_input_r[115];
assign temp_mult[116] = 16'd1711 * d1_input_r[116];
assign temp_mult[117] = 16'd2660 * d1_input_r[117];
assign temp_mult[118] = 16'd33161 * d1_input_r[118];
assign temp_mult[119] = 16'd2370 * d1_input_r[119];
assign temp_mult[120] = 16'd458 * d1_input_r[120];
assign temp_mult[121] = 16'd33115 * d1_input_r[121];
assign temp_mult[122] = 16'd34893 * d1_input_r[122];
assign temp_mult[123] = 16'd33368 * d1_input_r[123];
assign temp_mult[124] = 16'd2285 * d1_input_r[124];
assign temp_mult[125] = 16'd415 * d1_input_r[125];
assign temp_mult[126] = 16'd656 * d1_input_r[126];
assign temp_mult[127] = 16'd147 * d1_input_r[127];
assign temp_mult[128] = 16'd1024 * d1_input_r[128];
assign temp_mult[129] = 16'd1619 * d1_input_r[129];
assign temp_mult[130] = 16'd1585 * d1_input_r[130];
assign temp_mult[131] = 16'd33496 * d1_input_r[131];
assign temp_mult[132] = 16'd34669 * d1_input_r[132];
assign temp_mult[133] = 16'd35444 * d1_input_r[133];
assign temp_mult[134] = 16'd34470 * d1_input_r[134];
assign temp_mult[135] = 16'd33334 * d1_input_r[135];
assign temp_mult[136] = 16'd2565 * d1_input_r[136];
assign temp_mult[137] = 16'd33420 * d1_input_r[137];
assign temp_mult[138] = 16'd35502 * d1_input_r[138];
assign temp_mult[139] = 16'd33781 * d1_input_r[139];
assign temp_mult[140] = 16'd2085 * d1_input_r[140];
assign temp_mult[141] = 16'd328 * d1_input_r[141];
assign temp_mult[142] = 16'd32903 * d1_input_r[142];
assign temp_mult[143] = 16'd33928 * d1_input_r[143];
assign temp_mult[144] = 16'd34128 * d1_input_r[144];
assign temp_mult[145] = 16'd34319 * d1_input_r[145];
assign temp_mult[146] = 16'd33171 * d1_input_r[146];
assign temp_mult[147] = 16'd34067 * d1_input_r[147];
assign temp_mult[148] = 16'd381 * d1_input_r[148];
assign temp_mult[149] = 16'd1803 * d1_input_r[149];
assign temp_mult[150] = 16'd110 * d1_input_r[150];
assign temp_mult[151] = 16'd33524 * d1_input_r[151];
assign temp_mult[152] = 16'd33441 * d1_input_r[152];
assign temp_mult[153] = 16'd1502 * d1_input_r[153];
assign temp_mult[154] = 16'd1843 * d1_input_r[154];
assign temp_mult[155] = 16'd33835 * d1_input_r[155];
assign temp_mult[156] = 16'd1056 * d1_input_r[156];
assign temp_mult[157] = 16'd573 * d1_input_r[157];
assign temp_mult[158] = 16'd33310 * d1_input_r[158];
assign temp_mult[159] = 16'd34185 * d1_input_r[159];
assign temp_mult[160] = 16'd378 * d1_input_r[160];
assign temp_mult[161] = 16'd32980 * d1_input_r[161];
assign temp_mult[162] = 16'd318 * d1_input_r[162];
assign temp_mult[163] = 16'd34115 * d1_input_r[163];
assign temp_mult[164] = 16'd740 * d1_input_r[164];
assign temp_mult[165] = 16'd33599 * d1_input_r[165];
assign temp_mult[166] = 16'd34725 * d1_input_r[166];
assign temp_mult[167] = 16'd555 * d1_input_r[167];
assign temp_mult[168] = 16'd33489 * d1_input_r[168];
assign temp_mult[169] = 16'd32988 * d1_input_r[169];
assign temp_mult[170] = 16'd136 * d1_input_r[170];
assign temp_mult[171] = 16'd33689 * d1_input_r[171];
assign temp_mult[172] = 16'd32816 * d1_input_r[172];
assign temp_mult[173] = 16'd1937 * d1_input_r[173];
assign temp_mult[174] = 16'd33731 * d1_input_r[174];
assign temp_mult[175] = 16'd1016 * d1_input_r[175];
assign temp_mult[176] = 16'd1585 * d1_input_r[176];
assign temp_mult[177] = 16'd462 * d1_input_r[177];
assign temp_mult[178] = 16'd33246 * d1_input_r[178];
assign temp_mult[179] = 16'd659 * d1_input_r[179];
assign temp_mult[180] = 16'd35100 * d1_input_r[180];
assign temp_mult[181] = 16'd33522 * d1_input_r[181];
assign temp_mult[182] = 16'd781 * d1_input_r[182];
assign temp_mult[183] = 16'd630 * d1_input_r[183];
assign temp_mult[184] = 16'd32788 * d1_input_r[184];
assign temp_mult[185] = 16'd33054 * d1_input_r[185];
assign temp_mult[186] = 16'd2849 * d1_input_r[186];
assign temp_mult[187] = 16'd2577 * d1_input_r[187];
assign temp_mult[188] = 16'd33140 * d1_input_r[188];
assign temp_mult[189] = 16'd1847 * d1_input_r[189];
assign temp_mult[190] = 16'd33543 * d1_input_r[190];
assign temp_mult[191] = 16'd1058 * d1_input_r[191];
assign temp_mult[192] = 16'd61 * d1_input_r[192];
assign temp_mult[193] = 16'd432 * d1_input_r[193];
assign temp_mult[194] = 16'd33782 * d1_input_r[194];
assign temp_mult[195] = 16'd33483 * d1_input_r[195];
assign temp_mult[196] = 16'd1453 * d1_input_r[196];
assign temp_mult[197] = 16'd1136 * d1_input_r[197];
assign temp_mult[198] = 16'd34849 * d1_input_r[198];
assign temp_mult[199] = 16'd2280 * d1_input_r[199];
assign temp_mult[200] = 16'd2566 * d1_input_r[200];
assign temp_mult[201] = 16'd34460 * d1_input_r[201];
assign temp_mult[202] = 16'd34294 * d1_input_r[202];
assign temp_mult[203] = 16'd1276 * d1_input_r[203];
assign temp_mult[204] = 16'd1970 * d1_input_r[204];
assign temp_mult[205] = 16'd34243 * d1_input_r[205];
assign temp_mult[206] = 16'd1322 * d1_input_r[206];
assign temp_mult[207] = 16'd34864 * d1_input_r[207];
assign temp_mult[208] = 16'd33303 * d1_input_r[208];
assign temp_mult[209] = 16'd407 * d1_input_r[209];
assign temp_mult[210] = 16'd1732 * d1_input_r[210];
assign temp_mult[211] = 16'd340 * d1_input_r[211];
assign temp_mult[212] = 16'd1022 * d1_input_r[212];
assign temp_mult[213] = 16'd34272 * d1_input_r[213];
assign temp_mult[214] = 16'd33965 * d1_input_r[214];
assign temp_mult[215] = 16'd1057 * d1_input_r[215];
assign temp_mult[216] = 16'd215 * d1_input_r[216];
assign temp_mult[217] = 16'd1738 * d1_input_r[217];
assign temp_mult[218] = 16'd1293 * d1_input_r[218];
assign temp_mult[219] = 16'd3146 * d1_input_r[219];
assign temp_mult[220] = 16'd1060 * d1_input_r[220];
assign temp_mult[221] = 16'd1543 * d1_input_r[221];
assign temp_mult[222] = 16'd296 * d1_input_r[222];
assign temp_mult[223] = 16'd33327 * d1_input_r[223];
assign temp_mult[224] = 16'd34496 * d1_input_r[224];
assign temp_mult[225] = 16'd33170 * d1_input_r[225];
assign temp_mult[226] = 16'd507 * d1_input_r[226];
assign temp_mult[227] = 16'd2815 * d1_input_r[227];
assign temp_mult[228] = 16'd33973 * d1_input_r[228];
assign temp_mult[229] = 16'd33730 * d1_input_r[229];
assign temp_mult[230] = 16'd33450 * d1_input_r[230];
assign temp_mult[231] = 16'd687 * d1_input_r[231];
assign temp_mult[232] = 16'd2561 * d1_input_r[232];
assign temp_mult[233] = 16'd34430 * d1_input_r[233];
assign temp_mult[234] = 16'd802 * d1_input_r[234];
assign temp_mult[235] = 16'd34961 * d1_input_r[235];
assign temp_mult[236] = 16'd1664 * d1_input_r[236];
assign temp_mult[237] = 16'd1431 * d1_input_r[237];
assign temp_mult[238] = 16'd799 * d1_input_r[238];
assign temp_mult[239] = 16'd34597 * d1_input_r[239];
assign temp_mult[240] = 16'd35550 * d1_input_r[240];
assign temp_mult[241] = 16'd831 * d1_input_r[241];
assign temp_mult[242] = 16'd717 * d1_input_r[242];
assign temp_mult[243] = 16'd33328 * d1_input_r[243];
assign temp_mult[244] = 16'd35745 * d1_input_r[244];
assign temp_mult[245] = 16'd33702 * d1_input_r[245];
assign temp_mult[246] = 16'd632 * d1_input_r[246];
assign temp_mult[247] = 16'd34382 * d1_input_r[247];
assign temp_mult[248] = 16'd520 * d1_input_r[248];
assign temp_mult[249] = 16'd1811 * d1_input_r[249];
assign temp_mult[250] = 16'd33937 * d1_input_r[250];
assign temp_mult[251] = 16'd2222 * d1_input_r[251];
assign temp_mult[252] = 16'd1776 * d1_input_r[252];
assign temp_mult[253] = 16'd862 * d1_input_r[253];
assign temp_mult[254] = 16'd34076 * d1_input_r[254];
assign temp_mult[255] = 16'd2403 * d1_input_r[255];
assign temp_mult[256] = 16'd1741 * d1_input_r[0];
assign temp_mult[257] = 16'd580 * d1_input_r[1];
assign temp_mult[258] = 16'd644 * d1_input_r[2];
assign temp_mult[259] = 16'd33412 * d1_input_r[3];
assign temp_mult[260] = 16'd33545 * d1_input_r[4];
assign temp_mult[261] = 16'd35146 * d1_input_r[5];
assign temp_mult[262] = 16'd1832 * d1_input_r[6];
assign temp_mult[263] = 16'd1903 * d1_input_r[7];
assign temp_mult[264] = 16'd1961 * d1_input_r[8];
assign temp_mult[265] = 16'd34914 * d1_input_r[9];
assign temp_mult[266] = 16'd2360 * d1_input_r[10];
assign temp_mult[267] = 16'd907 * d1_input_r[11];
assign temp_mult[268] = 16'd32869 * d1_input_r[12];
assign temp_mult[269] = 16'd33679 * d1_input_r[13];
assign temp_mult[270] = 16'd32944 * d1_input_r[14];
assign temp_mult[271] = 16'd600 * d1_input_r[15];
assign temp_mult[272] = 16'd1603 * d1_input_r[16];
assign temp_mult[273] = 16'd33544 * d1_input_r[17];
assign temp_mult[274] = 16'd35058 * d1_input_r[18];
assign temp_mult[275] = 16'd32895 * d1_input_r[19];
assign temp_mult[276] = 16'd33413 * d1_input_r[20];
assign temp_mult[277] = 16'd35193 * d1_input_r[21];
assign temp_mult[278] = 16'd858 * d1_input_r[22];
assign temp_mult[279] = 16'd1606 * d1_input_r[23];
assign temp_mult[280] = 16'd1359 * d1_input_r[24];
assign temp_mult[281] = 16'd359 * d1_input_r[25];
assign temp_mult[282] = 16'd1545 * d1_input_r[26];
assign temp_mult[283] = 16'd33911 * d1_input_r[27];
assign temp_mult[284] = 16'd132 * d1_input_r[28];
assign temp_mult[285] = 16'd35108 * d1_input_r[29];
assign temp_mult[286] = 16'd34614 * d1_input_r[30];
assign temp_mult[287] = 16'd33613 * d1_input_r[31];
assign temp_mult[288] = 16'd33508 * d1_input_r[32];
assign temp_mult[289] = 16'd1699 * d1_input_r[33];
assign temp_mult[290] = 16'd34507 * d1_input_r[34];
assign temp_mult[291] = 16'd2576 * d1_input_r[35];
assign temp_mult[292] = 16'd994 * d1_input_r[36];
assign temp_mult[293] = 16'd178 * d1_input_r[37];
assign temp_mult[294] = 16'd32786 * d1_input_r[38];
assign temp_mult[295] = 16'd33136 * d1_input_r[39];
assign temp_mult[296] = 16'd2550 * d1_input_r[40];
assign temp_mult[297] = 16'd34846 * d1_input_r[41];
assign temp_mult[298] = 16'd33587 * d1_input_r[42];
assign temp_mult[299] = 16'd34555 * d1_input_r[43];
assign temp_mult[300] = 16'd35646 * d1_input_r[44];
assign temp_mult[301] = 16'd34822 * d1_input_r[45];
assign temp_mult[302] = 16'd866 * d1_input_r[46];
assign temp_mult[303] = 16'd33467 * d1_input_r[47];
assign temp_mult[304] = 16'd1925 * d1_input_r[48];
assign temp_mult[305] = 16'd532 * d1_input_r[49];
assign temp_mult[306] = 16'd1213 * d1_input_r[50];
assign temp_mult[307] = 16'd1065 * d1_input_r[51];
assign temp_mult[308] = 16'd34078 * d1_input_r[52];
assign temp_mult[309] = 16'd33242 * d1_input_r[53];
assign temp_mult[310] = 16'd1949 * d1_input_r[54];
assign temp_mult[311] = 16'd33600 * d1_input_r[55];
assign temp_mult[312] = 16'd915 * d1_input_r[56];
assign temp_mult[313] = 16'd1177 * d1_input_r[57];
assign temp_mult[314] = 16'd34051 * d1_input_r[58];
assign temp_mult[315] = 16'd1066 * d1_input_r[59];
assign temp_mult[316] = 16'd1121 * d1_input_r[60];
assign temp_mult[317] = 16'd33143 * d1_input_r[61];
assign temp_mult[318] = 16'd34049 * d1_input_r[62];
assign temp_mult[319] = 16'd1024 * d1_input_r[63];
assign temp_mult[320] = 16'd449 * d1_input_r[64];
assign temp_mult[321] = 16'd34668 * d1_input_r[65];
assign temp_mult[322] = 16'd175 * d1_input_r[66];
assign temp_mult[323] = 16'd34370 * d1_input_r[67];
assign temp_mult[324] = 16'd131 * d1_input_r[68];
assign temp_mult[325] = 16'd34900 * d1_input_r[69];
assign temp_mult[326] = 16'd169 * d1_input_r[70];
assign temp_mult[327] = 16'd1022 * d1_input_r[71];
assign temp_mult[328] = 16'd767 * d1_input_r[72];
assign temp_mult[329] = 16'd35378 * d1_input_r[73];
assign temp_mult[330] = 16'd106 * d1_input_r[74];
assign temp_mult[331] = 16'd964 * d1_input_r[75];
assign temp_mult[332] = 16'd33114 * d1_input_r[76];
assign temp_mult[333] = 16'd407 * d1_input_r[77];
assign temp_mult[334] = 16'd1887 * d1_input_r[78];
assign temp_mult[335] = 16'd35161 * d1_input_r[79];
assign temp_mult[336] = 16'd34277 * d1_input_r[80];
assign temp_mult[337] = 16'd962 * d1_input_r[81];
assign temp_mult[338] = 16'd1023 * d1_input_r[82];
assign temp_mult[339] = 16'd35844 * d1_input_r[83];
assign temp_mult[340] = 16'd1524 * d1_input_r[84];
assign temp_mult[341] = 16'd3028 * d1_input_r[85];
assign temp_mult[342] = 16'd33678 * d1_input_r[86];
assign temp_mult[343] = 16'd33406 * d1_input_r[87];
assign temp_mult[344] = 16'd1591 * d1_input_r[88];
assign temp_mult[345] = 16'd1445 * d1_input_r[89];
assign temp_mult[346] = 16'd34257 * d1_input_r[90];
assign temp_mult[347] = 16'd33017 * d1_input_r[91];
assign temp_mult[348] = 16'd184 * d1_input_r[92];
assign temp_mult[349] = 16'd811 * d1_input_r[93];
assign temp_mult[350] = 16'd34839 * d1_input_r[94];
assign temp_mult[351] = 16'd2238 * d1_input_r[95];
assign temp_mult[352] = 16'd34491 * d1_input_r[96];
assign temp_mult[353] = 16'd579 * d1_input_r[97];
assign temp_mult[354] = 16'd1670 * d1_input_r[98];
assign temp_mult[355] = 16'd1554 * d1_input_r[99];
assign temp_mult[356] = 16'd34742 * d1_input_r[100];
assign temp_mult[357] = 16'd1031 * d1_input_r[101];
assign temp_mult[358] = 16'd1224 * d1_input_r[102];
assign temp_mult[359] = 16'd2158 * d1_input_r[103];
assign temp_mult[360] = 16'd1880 * d1_input_r[104];
assign temp_mult[361] = 16'd32913 * d1_input_r[105];
assign temp_mult[362] = 16'd33427 * d1_input_r[106];
assign temp_mult[363] = 16'd2340 * d1_input_r[107];
assign temp_mult[364] = 16'd34072 * d1_input_r[108];
assign temp_mult[365] = 16'd32983 * d1_input_r[109];
assign temp_mult[366] = 16'd34055 * d1_input_r[110];
assign temp_mult[367] = 16'd544 * d1_input_r[111];
assign temp_mult[368] = 16'd34468 * d1_input_r[112];
assign temp_mult[369] = 16'd2794 * d1_input_r[113];
assign temp_mult[370] = 16'd32841 * d1_input_r[114];
assign temp_mult[371] = 16'd33397 * d1_input_r[115];
assign temp_mult[372] = 16'd605 * d1_input_r[116];
assign temp_mult[373] = 16'd33916 * d1_input_r[117];
assign temp_mult[374] = 16'd33556 * d1_input_r[118];
assign temp_mult[375] = 16'd34927 * d1_input_r[119];
assign temp_mult[376] = 16'd580 * d1_input_r[120];
assign temp_mult[377] = 16'd1346 * d1_input_r[121];
assign temp_mult[378] = 16'd530 * d1_input_r[122];
assign temp_mult[379] = 16'd33930 * d1_input_r[123];
assign temp_mult[380] = 16'd1364 * d1_input_r[124];
assign temp_mult[381] = 16'd1351 * d1_input_r[125];
assign temp_mult[382] = 16'd2027 * d1_input_r[126];
assign temp_mult[383] = 16'd33636 * d1_input_r[127];
assign temp_mult[384] = 16'd420 * d1_input_r[128];
assign temp_mult[385] = 16'd35008 * d1_input_r[129];
assign temp_mult[386] = 16'd34166 * d1_input_r[130];
assign temp_mult[387] = 16'd33450 * d1_input_r[131];
assign temp_mult[388] = 16'd34803 * d1_input_r[132];
assign temp_mult[389] = 16'd35081 * d1_input_r[133];
assign temp_mult[390] = 16'd35312 * d1_input_r[134];
assign temp_mult[391] = 16'd3088 * d1_input_r[135];
assign temp_mult[392] = 16'd2911 * d1_input_r[136];
assign temp_mult[393] = 16'd1473 * d1_input_r[137];
assign temp_mult[394] = 16'd1851 * d1_input_r[138];
assign temp_mult[395] = 16'd752 * d1_input_r[139];
assign temp_mult[396] = 16'd33051 * d1_input_r[140];
assign temp_mult[397] = 16'd2588 * d1_input_r[141];
assign temp_mult[398] = 16'd9 * d1_input_r[142];
assign temp_mult[399] = 16'd919 * d1_input_r[143];
assign temp_mult[400] = 16'd82 * d1_input_r[144];
assign temp_mult[401] = 16'd1822 * d1_input_r[145];
assign temp_mult[402] = 16'd33799 * d1_input_r[146];
assign temp_mult[403] = 16'd35337 * d1_input_r[147];
assign temp_mult[404] = 16'd1641 * d1_input_r[148];
assign temp_mult[405] = 16'd34106 * d1_input_r[149];
assign temp_mult[406] = 16'd33158 * d1_input_r[150];
assign temp_mult[407] = 16'd534 * d1_input_r[151];
assign temp_mult[408] = 16'd1553 * d1_input_r[152];
assign temp_mult[409] = 16'd35250 * d1_input_r[153];
assign temp_mult[410] = 16'd552 * d1_input_r[154];
assign temp_mult[411] = 16'd1387 * d1_input_r[155];
assign temp_mult[412] = 16'd2896 * d1_input_r[156];
assign temp_mult[413] = 16'd33531 * d1_input_r[157];
assign temp_mult[414] = 16'd34582 * d1_input_r[158];
assign temp_mult[415] = 16'd590 * d1_input_r[159];
assign temp_mult[416] = 16'd34816 * d1_input_r[160];
assign temp_mult[417] = 16'd34292 * d1_input_r[161];
assign temp_mult[418] = 16'd90 * d1_input_r[162];
assign temp_mult[419] = 16'd1120 * d1_input_r[163];
assign temp_mult[420] = 16'd416 * d1_input_r[164];
assign temp_mult[421] = 16'd34664 * d1_input_r[165];
assign temp_mult[422] = 16'd543 * d1_input_r[166];
assign temp_mult[423] = 16'd2847 * d1_input_r[167];
assign temp_mult[424] = 16'd1904 * d1_input_r[168];
assign temp_mult[425] = 16'd34336 * d1_input_r[169];
assign temp_mult[426] = 16'd34073 * d1_input_r[170];
assign temp_mult[427] = 16'd33829 * d1_input_r[171];
assign temp_mult[428] = 16'd13 * d1_input_r[172];
assign temp_mult[429] = 16'd454 * d1_input_r[173];
assign temp_mult[430] = 16'd34606 * d1_input_r[174];
assign temp_mult[431] = 16'd32777 * d1_input_r[175];
assign temp_mult[432] = 16'd150 * d1_input_r[176];
assign temp_mult[433] = 16'd32839 * d1_input_r[177];
assign temp_mult[434] = 16'd1999 * d1_input_r[178];
assign temp_mult[435] = 16'd34879 * d1_input_r[179];
assign temp_mult[436] = 16'd63 * d1_input_r[180];
assign temp_mult[437] = 16'd33351 * d1_input_r[181];
assign temp_mult[438] = 16'd393 * d1_input_r[182];
assign temp_mult[439] = 16'd33995 * d1_input_r[183];
assign temp_mult[440] = 16'd895 * d1_input_r[184];
assign temp_mult[441] = 16'd1694 * d1_input_r[185];
assign temp_mult[442] = 16'd248 * d1_input_r[186];
assign temp_mult[443] = 16'd33020 * d1_input_r[187];
assign temp_mult[444] = 16'd32832 * d1_input_r[188];
assign temp_mult[445] = 16'd33787 * d1_input_r[189];
assign temp_mult[446] = 16'd35556 * d1_input_r[190];
assign temp_mult[447] = 16'd32810 * d1_input_r[191];
assign temp_mult[448] = 16'd34013 * d1_input_r[192];
assign temp_mult[449] = 16'd32872 * d1_input_r[193];
assign temp_mult[450] = 16'd34942 * d1_input_r[194];
assign temp_mult[451] = 16'd2430 * d1_input_r[195];
assign temp_mult[452] = 16'd3005 * d1_input_r[196];
assign temp_mult[453] = 16'd1292 * d1_input_r[197];
assign temp_mult[454] = 16'd480 * d1_input_r[198];
assign temp_mult[455] = 16'd33888 * d1_input_r[199];
assign temp_mult[456] = 16'd149 * d1_input_r[200];
assign temp_mult[457] = 16'd33879 * d1_input_r[201];
assign temp_mult[458] = 16'd776 * d1_input_r[202];
assign temp_mult[459] = 16'd34760 * d1_input_r[203];
assign temp_mult[460] = 16'd545 * d1_input_r[204];
assign temp_mult[461] = 16'd33914 * d1_input_r[205];
assign temp_mult[462] = 16'd34264 * d1_input_r[206];
assign temp_mult[463] = 16'd32956 * d1_input_r[207];
assign temp_mult[464] = 16'd35715 * d1_input_r[208];
assign temp_mult[465] = 16'd33075 * d1_input_r[209];
assign temp_mult[466] = 16'd1946 * d1_input_r[210];
assign temp_mult[467] = 16'd2275 * d1_input_r[211];
assign temp_mult[468] = 16'd239 * d1_input_r[212];
assign temp_mult[469] = 16'd35785 * d1_input_r[213];
assign temp_mult[470] = 16'd33729 * d1_input_r[214];
assign temp_mult[471] = 16'd691 * d1_input_r[215];
assign temp_mult[472] = 16'd1719 * d1_input_r[216];
assign temp_mult[473] = 16'd34842 * d1_input_r[217];
assign temp_mult[474] = 16'd33631 * d1_input_r[218];
assign temp_mult[475] = 16'd2998 * d1_input_r[219];
assign temp_mult[476] = 16'd73 * d1_input_r[220];
assign temp_mult[477] = 16'd1222 * d1_input_r[221];
assign temp_mult[478] = 16'd35619 * d1_input_r[222];
assign temp_mult[479] = 16'd1577 * d1_input_r[223];
assign temp_mult[480] = 16'd327 * d1_input_r[224];
assign temp_mult[481] = 16'd921 * d1_input_r[225];
assign temp_mult[482] = 16'd33839 * d1_input_r[226];
assign temp_mult[483] = 16'd2244 * d1_input_r[227];
assign temp_mult[484] = 16'd33637 * d1_input_r[228];
assign temp_mult[485] = 16'd33625 * d1_input_r[229];
assign temp_mult[486] = 16'd1644 * d1_input_r[230];
assign temp_mult[487] = 16'd33886 * d1_input_r[231];
assign temp_mult[488] = 16'd34508 * d1_input_r[232];
assign temp_mult[489] = 16'd33641 * d1_input_r[233];
assign temp_mult[490] = 16'd678 * d1_input_r[234];
assign temp_mult[491] = 16'd1838 * d1_input_r[235];
assign temp_mult[492] = 16'd34908 * d1_input_r[236];
assign temp_mult[493] = 16'd2054 * d1_input_r[237];
assign temp_mult[494] = 16'd802 * d1_input_r[238];
assign temp_mult[495] = 16'd34375 * d1_input_r[239];
assign temp_mult[496] = 16'd1084 * d1_input_r[240];
assign temp_mult[497] = 16'd1963 * d1_input_r[241];
assign temp_mult[498] = 16'd34540 * d1_input_r[242];
assign temp_mult[499] = 16'd1779 * d1_input_r[243];
assign temp_mult[500] = 16'd33956 * d1_input_r[244];
assign temp_mult[501] = 16'd33525 * d1_input_r[245];
assign temp_mult[502] = 16'd208 * d1_input_r[246];
assign temp_mult[503] = 16'd32888 * d1_input_r[247];
assign temp_mult[504] = 16'd1170 * d1_input_r[248];
assign temp_mult[505] = 16'd35266 * d1_input_r[249];
assign temp_mult[506] = 16'd620 * d1_input_r[250];
assign temp_mult[507] = 16'd344 * d1_input_r[251];
assign temp_mult[508] = 16'd1267 * d1_input_r[252];
assign temp_mult[509] = 16'd1764 * d1_input_r[253];
assign temp_mult[510] = 16'd33316 * d1_input_r[254];
assign temp_mult[511] = 16'd34 * d1_input_r[255];
assign temp_mult[512] = 16'd34854 * d1_input_r[0];
assign temp_mult[513] = 16'd32894 * d1_input_r[1];
assign temp_mult[514] = 16'd33087 * d1_input_r[2];
assign temp_mult[515] = 16'd35780 * d1_input_r[3];
assign temp_mult[516] = 16'd32938 * d1_input_r[4];
assign temp_mult[517] = 16'd3115 * d1_input_r[5];
assign temp_mult[518] = 16'd33788 * d1_input_r[6];
assign temp_mult[519] = 16'd1665 * d1_input_r[7];
assign temp_mult[520] = 16'd255 * d1_input_r[8];
assign temp_mult[521] = 16'd33302 * d1_input_r[9];
assign temp_mult[522] = 16'd35635 * d1_input_r[10];
assign temp_mult[523] = 16'd1048 * d1_input_r[11];
assign temp_mult[524] = 16'd32993 * d1_input_r[12];
assign temp_mult[525] = 16'd33350 * d1_input_r[13];
assign temp_mult[526] = 16'd34291 * d1_input_r[14];
assign temp_mult[527] = 16'd34515 * d1_input_r[15];
assign temp_mult[528] = 16'd2179 * d1_input_r[16];
assign temp_mult[529] = 16'd150 * d1_input_r[17];
assign temp_mult[530] = 16'd2025 * d1_input_r[18];
assign temp_mult[531] = 16'd33532 * d1_input_r[19];
assign temp_mult[532] = 16'd33189 * d1_input_r[20];
assign temp_mult[533] = 16'd1410 * d1_input_r[21];
assign temp_mult[534] = 16'd548 * d1_input_r[22];
assign temp_mult[535] = 16'd36 * d1_input_r[23];
assign temp_mult[536] = 16'd33979 * d1_input_r[24];
assign temp_mult[537] = 16'd878 * d1_input_r[25];
assign temp_mult[538] = 16'd2624 * d1_input_r[26];
assign temp_mult[539] = 16'd964 * d1_input_r[27];
assign temp_mult[540] = 16'd1693 * d1_input_r[28];
assign temp_mult[541] = 16'd906 * d1_input_r[29];
assign temp_mult[542] = 16'd1792 * d1_input_r[30];
assign temp_mult[543] = 16'd35761 * d1_input_r[31];
assign temp_mult[544] = 16'd33414 * d1_input_r[32];
assign temp_mult[545] = 16'd1335 * d1_input_r[33];
assign temp_mult[546] = 16'd34930 * d1_input_r[34];
assign temp_mult[547] = 16'd34174 * d1_input_r[35];
assign temp_mult[548] = 16'd1260 * d1_input_r[36];
assign temp_mult[549] = 16'd33425 * d1_input_r[37];
assign temp_mult[550] = 16'd35336 * d1_input_r[38];
assign temp_mult[551] = 16'd1229 * d1_input_r[39];
assign temp_mult[552] = 16'd1304 * d1_input_r[40];
assign temp_mult[553] = 16'd196 * d1_input_r[41];
assign temp_mult[554] = 16'd506 * d1_input_r[42];
assign temp_mult[555] = 16'd35113 * d1_input_r[43];
assign temp_mult[556] = 16'd2856 * d1_input_r[44];
assign temp_mult[557] = 16'd1360 * d1_input_r[45];
assign temp_mult[558] = 16'd34558 * d1_input_r[46];
assign temp_mult[559] = 16'd34245 * d1_input_r[47];
assign temp_mult[560] = 16'd829 * d1_input_r[48];
assign temp_mult[561] = 16'd126 * d1_input_r[49];
assign temp_mult[562] = 16'd32871 * d1_input_r[50];
assign temp_mult[563] = 16'd118 * d1_input_r[51];
assign temp_mult[564] = 16'd33735 * d1_input_r[52];
assign temp_mult[565] = 16'd34828 * d1_input_r[53];
assign temp_mult[566] = 16'd33243 * d1_input_r[54];
assign temp_mult[567] = 16'd2425 * d1_input_r[55];
assign temp_mult[568] = 16'd35539 * d1_input_r[56];
assign temp_mult[569] = 16'd34095 * d1_input_r[57];
assign temp_mult[570] = 16'd33530 * d1_input_r[58];
assign temp_mult[571] = 16'd34354 * d1_input_r[59];
assign temp_mult[572] = 16'd33064 * d1_input_r[60];
assign temp_mult[573] = 16'd1119 * d1_input_r[61];
assign temp_mult[574] = 16'd34288 * d1_input_r[62];
assign temp_mult[575] = 16'd754 * d1_input_r[63];
assign temp_mult[576] = 16'd33814 * d1_input_r[64];
assign temp_mult[577] = 16'd33496 * d1_input_r[65];
assign temp_mult[578] = 16'd1002 * d1_input_r[66];
assign temp_mult[579] = 16'd35658 * d1_input_r[67];
assign temp_mult[580] = 16'd34031 * d1_input_r[68];
assign temp_mult[581] = 16'd2293 * d1_input_r[69];
assign temp_mult[582] = 16'd1847 * d1_input_r[70];
assign temp_mult[583] = 16'd34447 * d1_input_r[71];
assign temp_mult[584] = 16'd34904 * d1_input_r[72];
assign temp_mult[585] = 16'd1708 * d1_input_r[73];
assign temp_mult[586] = 16'd33147 * d1_input_r[74];
assign temp_mult[587] = 16'd814 * d1_input_r[75];
assign temp_mult[588] = 16'd2926 * d1_input_r[76];
assign temp_mult[589] = 16'd2192 * d1_input_r[77];
assign temp_mult[590] = 16'd689 * d1_input_r[78];
assign temp_mult[591] = 16'd33769 * d1_input_r[79];
assign temp_mult[592] = 16'd33866 * d1_input_r[80];
assign temp_mult[593] = 16'd34800 * d1_input_r[81];
assign temp_mult[594] = 16'd33957 * d1_input_r[82];
assign temp_mult[595] = 16'd2888 * d1_input_r[83];
assign temp_mult[596] = 16'd34461 * d1_input_r[84];
assign temp_mult[597] = 16'd35748 * d1_input_r[85];
assign temp_mult[598] = 16'd1750 * d1_input_r[86];
assign temp_mult[599] = 16'd32950 * d1_input_r[87];
assign temp_mult[600] = 16'd35135 * d1_input_r[88];
assign temp_mult[601] = 16'd600 * d1_input_r[89];
assign temp_mult[602] = 16'd1379 * d1_input_r[90];
assign temp_mult[603] = 16'd35741 * d1_input_r[91];
assign temp_mult[604] = 16'd34353 * d1_input_r[92];
assign temp_mult[605] = 16'd2396 * d1_input_r[93];
assign temp_mult[606] = 16'd859 * d1_input_r[94];
assign temp_mult[607] = 16'd34582 * d1_input_r[95];
assign temp_mult[608] = 16'd646 * d1_input_r[96];
assign temp_mult[609] = 16'd1326 * d1_input_r[97];
assign temp_mult[610] = 16'd35144 * d1_input_r[98];
assign temp_mult[611] = 16'd33240 * d1_input_r[99];
assign temp_mult[612] = 16'd33956 * d1_input_r[100];
assign temp_mult[613] = 16'd32832 * d1_input_r[101];
assign temp_mult[614] = 16'd34316 * d1_input_r[102];
assign temp_mult[615] = 16'd698 * d1_input_r[103];
assign temp_mult[616] = 16'd1393 * d1_input_r[104];
assign temp_mult[617] = 16'd1141 * d1_input_r[105];
assign temp_mult[618] = 16'd972 * d1_input_r[106];
assign temp_mult[619] = 16'd34911 * d1_input_r[107];
assign temp_mult[620] = 16'd32945 * d1_input_r[108];
assign temp_mult[621] = 16'd1092 * d1_input_r[109];
assign temp_mult[622] = 16'd33433 * d1_input_r[110];
assign temp_mult[623] = 16'd33893 * d1_input_r[111];
assign temp_mult[624] = 16'd32849 * d1_input_r[112];
assign temp_mult[625] = 16'd35215 * d1_input_r[113];
assign temp_mult[626] = 16'd34464 * d1_input_r[114];
assign temp_mult[627] = 16'd1878 * d1_input_r[115];
assign temp_mult[628] = 16'd33327 * d1_input_r[116];
assign temp_mult[629] = 16'd722 * d1_input_r[117];
assign temp_mult[630] = 16'd35433 * d1_input_r[118];
assign temp_mult[631] = 16'd791 * d1_input_r[119];
assign temp_mult[632] = 16'd100 * d1_input_r[120];
assign temp_mult[633] = 16'd34389 * d1_input_r[121];
assign temp_mult[634] = 16'd33590 * d1_input_r[122];
assign temp_mult[635] = 16'd35287 * d1_input_r[123];
assign temp_mult[636] = 16'd35240 * d1_input_r[124];
assign temp_mult[637] = 16'd1563 * d1_input_r[125];
assign temp_mult[638] = 16'd34498 * d1_input_r[126];
assign temp_mult[639] = 16'd35617 * d1_input_r[127];
assign temp_mult[640] = 16'd33841 * d1_input_r[128];
assign temp_mult[641] = 16'd1287 * d1_input_r[129];
assign temp_mult[642] = 16'd1636 * d1_input_r[130];
assign temp_mult[643] = 16'd34680 * d1_input_r[131];
assign temp_mult[644] = 16'd1541 * d1_input_r[132];
assign temp_mult[645] = 16'd1766 * d1_input_r[133];
assign temp_mult[646] = 16'd1920 * d1_input_r[134];
assign temp_mult[647] = 16'd35818 * d1_input_r[135];
assign temp_mult[648] = 16'd1451 * d1_input_r[136];
assign temp_mult[649] = 16'd2417 * d1_input_r[137];
assign temp_mult[650] = 16'd34665 * d1_input_r[138];
assign temp_mult[651] = 16'd2462 * d1_input_r[139];
assign temp_mult[652] = 16'd33322 * d1_input_r[140];
assign temp_mult[653] = 16'd35852 * d1_input_r[141];
assign temp_mult[654] = 16'd33083 * d1_input_r[142];
assign temp_mult[655] = 16'd32940 * d1_input_r[143];
assign temp_mult[656] = 16'd1868 * d1_input_r[144];
assign temp_mult[657] = 16'd35512 * d1_input_r[145];
assign temp_mult[658] = 16'd33088 * d1_input_r[146];
assign temp_mult[659] = 16'd33373 * d1_input_r[147];
assign temp_mult[660] = 16'd32838 * d1_input_r[148];
assign temp_mult[661] = 16'd33159 * d1_input_r[149];
assign temp_mult[662] = 16'd225 * d1_input_r[150];
assign temp_mult[663] = 16'd1899 * d1_input_r[151];
assign temp_mult[664] = 16'd33463 * d1_input_r[152];
assign temp_mult[665] = 16'd264 * d1_input_r[153];
assign temp_mult[666] = 16'd33642 * d1_input_r[154];
assign temp_mult[667] = 16'd33501 * d1_input_r[155];
assign temp_mult[668] = 16'd1393 * d1_input_r[156];
assign temp_mult[669] = 16'd34539 * d1_input_r[157];
assign temp_mult[670] = 16'd32901 * d1_input_r[158];
assign temp_mult[671] = 16'd34254 * d1_input_r[159];
assign temp_mult[672] = 16'd33101 * d1_input_r[160];
assign temp_mult[673] = 16'd33289 * d1_input_r[161];
assign temp_mult[674] = 16'd34653 * d1_input_r[162];
assign temp_mult[675] = 16'd32795 * d1_input_r[163];
assign temp_mult[676] = 16'd35440 * d1_input_r[164];
assign temp_mult[677] = 16'd33852 * d1_input_r[165];
assign temp_mult[678] = 16'd756 * d1_input_r[166];
assign temp_mult[679] = 16'd35268 * d1_input_r[167];
assign temp_mult[680] = 16'd1808 * d1_input_r[168];
assign temp_mult[681] = 16'd33602 * d1_input_r[169];
assign temp_mult[682] = 16'd1456 * d1_input_r[170];
assign temp_mult[683] = 16'd32960 * d1_input_r[171];
assign temp_mult[684] = 16'd34305 * d1_input_r[172];
assign temp_mult[685] = 16'd955 * d1_input_r[173];
assign temp_mult[686] = 16'd32814 * d1_input_r[174];
assign temp_mult[687] = 16'd1790 * d1_input_r[175];
assign temp_mult[688] = 16'd404 * d1_input_r[176];
assign temp_mult[689] = 16'd33401 * d1_input_r[177];
assign temp_mult[690] = 16'd598 * d1_input_r[178];
assign temp_mult[691] = 16'd34933 * d1_input_r[179];
assign temp_mult[692] = 16'd34034 * d1_input_r[180];
assign temp_mult[693] = 16'd2652 * d1_input_r[181];
assign temp_mult[694] = 16'd1940 * d1_input_r[182];
assign temp_mult[695] = 16'd33622 * d1_input_r[183];
assign temp_mult[696] = 16'd34213 * d1_input_r[184];
assign temp_mult[697] = 16'd32877 * d1_input_r[185];
assign temp_mult[698] = 16'd34691 * d1_input_r[186];
assign temp_mult[699] = 16'd1503 * d1_input_r[187];
assign temp_mult[700] = 16'd1608 * d1_input_r[188];
assign temp_mult[701] = 16'd34270 * d1_input_r[189];
assign temp_mult[702] = 16'd508 * d1_input_r[190];
assign temp_mult[703] = 16'd35404 * d1_input_r[191];
assign temp_mult[704] = 16'd34417 * d1_input_r[192];
assign temp_mult[705] = 16'd973 * d1_input_r[193];
assign temp_mult[706] = 16'd35455 * d1_input_r[194];
assign temp_mult[707] = 16'd33200 * d1_input_r[195];
assign temp_mult[708] = 16'd34772 * d1_input_r[196];
assign temp_mult[709] = 16'd335 * d1_input_r[197];
assign temp_mult[710] = 16'd33776 * d1_input_r[198];
assign temp_mult[711] = 16'd1079 * d1_input_r[199];
assign temp_mult[712] = 16'd34333 * d1_input_r[200];
assign temp_mult[713] = 16'd33480 * d1_input_r[201];
assign temp_mult[714] = 16'd33876 * d1_input_r[202];
assign temp_mult[715] = 16'd110 * d1_input_r[203];
assign temp_mult[716] = 16'd35795 * d1_input_r[204];
assign temp_mult[717] = 16'd35338 * d1_input_r[205];
assign temp_mult[718] = 16'd34021 * d1_input_r[206];
assign temp_mult[719] = 16'd2448 * d1_input_r[207];
assign temp_mult[720] = 16'd2575 * d1_input_r[208];
assign temp_mult[721] = 16'd1248 * d1_input_r[209];
assign temp_mult[722] = 16'd1278 * d1_input_r[210];
assign temp_mult[723] = 16'd574 * d1_input_r[211];
assign temp_mult[724] = 16'd1197 * d1_input_r[212];
assign temp_mult[725] = 16'd2244 * d1_input_r[213];
assign temp_mult[726] = 16'd671 * d1_input_r[214];
assign temp_mult[727] = 16'd32774 * d1_input_r[215];
assign temp_mult[728] = 16'd883 * d1_input_r[216];
assign temp_mult[729] = 16'd914 * d1_input_r[217];
assign temp_mult[730] = 16'd35121 * d1_input_r[218];
assign temp_mult[731] = 16'd534 * d1_input_r[219];
assign temp_mult[732] = 16'd32856 * d1_input_r[220];
assign temp_mult[733] = 16'd33641 * d1_input_r[221];
assign temp_mult[734] = 16'd786 * d1_input_r[222];
assign temp_mult[735] = 16'd44 * d1_input_r[223];
assign temp_mult[736] = 16'd35437 * d1_input_r[224];
assign temp_mult[737] = 16'd1231 * d1_input_r[225];
assign temp_mult[738] = 16'd2247 * d1_input_r[226];
assign temp_mult[739] = 16'd1578 * d1_input_r[227];
assign temp_mult[740] = 16'd32935 * d1_input_r[228];
assign temp_mult[741] = 16'd33113 * d1_input_r[229];
assign temp_mult[742] = 16'd33153 * d1_input_r[230];
assign temp_mult[743] = 16'd1108 * d1_input_r[231];
assign temp_mult[744] = 16'd34843 * d1_input_r[232];
assign temp_mult[745] = 16'd625 * d1_input_r[233];
assign temp_mult[746] = 16'd2587 * d1_input_r[234];
assign temp_mult[747] = 16'd34189 * d1_input_r[235];
assign temp_mult[748] = 16'd2606 * d1_input_r[236];
assign temp_mult[749] = 16'd34205 * d1_input_r[237];
assign temp_mult[750] = 16'd33968 * d1_input_r[238];
assign temp_mult[751] = 16'd2741 * d1_input_r[239];
assign temp_mult[752] = 16'd1787 * d1_input_r[240];
assign temp_mult[753] = 16'd34089 * d1_input_r[241];
assign temp_mult[754] = 16'd33357 * d1_input_r[242];
assign temp_mult[755] = 16'd35082 * d1_input_r[243];
assign temp_mult[756] = 16'd413 * d1_input_r[244];
assign temp_mult[757] = 16'd34451 * d1_input_r[245];
assign temp_mult[758] = 16'd813 * d1_input_r[246];
assign temp_mult[759] = 16'd35048 * d1_input_r[247];
assign temp_mult[760] = 16'd34781 * d1_input_r[248];
assign temp_mult[761] = 16'd2325 * d1_input_r[249];
assign temp_mult[762] = 16'd32962 * d1_input_r[250];
assign temp_mult[763] = 16'd33548 * d1_input_r[251];
assign temp_mult[764] = 16'd728 * d1_input_r[252];
assign temp_mult[765] = 16'd1957 * d1_input_r[253];
assign temp_mult[766] = 16'd33473 * d1_input_r[254];
assign temp_mult[767] = 16'd35034 * d1_input_r[255];
assign temp_mult[768] = 16'd34438 * d1_input_r[0];
assign temp_mult[769] = 16'd341 * d1_input_r[1];
assign temp_mult[770] = 16'd2510 * d1_input_r[2];
assign temp_mult[771] = 16'd35385 * d1_input_r[3];
assign temp_mult[772] = 16'd33538 * d1_input_r[4];
assign temp_mult[773] = 16'd1219 * d1_input_r[5];
assign temp_mult[774] = 16'd34335 * d1_input_r[6];
assign temp_mult[775] = 16'd359 * d1_input_r[7];
assign temp_mult[776] = 16'd33769 * d1_input_r[8];
assign temp_mult[777] = 16'd785 * d1_input_r[9];
assign temp_mult[778] = 16'd795 * d1_input_r[10];
assign temp_mult[779] = 16'd34594 * d1_input_r[11];
assign temp_mult[780] = 16'd32802 * d1_input_r[12];
assign temp_mult[781] = 16'd218 * d1_input_r[13];
assign temp_mult[782] = 16'd35876 * d1_input_r[14];
assign temp_mult[783] = 16'd34609 * d1_input_r[15];
assign temp_mult[784] = 16'd33842 * d1_input_r[16];
assign temp_mult[785] = 16'd2030 * d1_input_r[17];
assign temp_mult[786] = 16'd1441 * d1_input_r[18];
assign temp_mult[787] = 16'd1348 * d1_input_r[19];
assign temp_mult[788] = 16'd2549 * d1_input_r[20];
assign temp_mult[789] = 16'd143 * d1_input_r[21];
assign temp_mult[790] = 16'd32903 * d1_input_r[22];
assign temp_mult[791] = 16'd893 * d1_input_r[23];
assign temp_mult[792] = 16'd33551 * d1_input_r[24];
assign temp_mult[793] = 16'd32940 * d1_input_r[25];
assign temp_mult[794] = 16'd33418 * d1_input_r[26];
assign temp_mult[795] = 16'd33002 * d1_input_r[27];
assign temp_mult[796] = 16'd1182 * d1_input_r[28];
assign temp_mult[797] = 16'd2320 * d1_input_r[29];
assign temp_mult[798] = 16'd33257 * d1_input_r[30];
assign temp_mult[799] = 16'd34917 * d1_input_r[31];
assign temp_mult[800] = 16'd34833 * d1_input_r[32];
assign temp_mult[801] = 16'd1530 * d1_input_r[33];
assign temp_mult[802] = 16'd33458 * d1_input_r[34];
assign temp_mult[803] = 16'd34845 * d1_input_r[35];
assign temp_mult[804] = 16'd34334 * d1_input_r[36];
assign temp_mult[805] = 16'd71 * d1_input_r[37];
assign temp_mult[806] = 16'd750 * d1_input_r[38];
assign temp_mult[807] = 16'd34882 * d1_input_r[39];
assign temp_mult[808] = 16'd315 * d1_input_r[40];
assign temp_mult[809] = 16'd34564 * d1_input_r[41];
assign temp_mult[810] = 16'd33520 * d1_input_r[42];
assign temp_mult[811] = 16'd34593 * d1_input_r[43];
assign temp_mult[812] = 16'd33381 * d1_input_r[44];
assign temp_mult[813] = 16'd1810 * d1_input_r[45];
assign temp_mult[814] = 16'd2352 * d1_input_r[46];
assign temp_mult[815] = 16'd2566 * d1_input_r[47];
assign temp_mult[816] = 16'd33629 * d1_input_r[48];
assign temp_mult[817] = 16'd420 * d1_input_r[49];
assign temp_mult[818] = 16'd2279 * d1_input_r[50];
assign temp_mult[819] = 16'd33448 * d1_input_r[51];
assign temp_mult[820] = 16'd34339 * d1_input_r[52];
assign temp_mult[821] = 16'd35377 * d1_input_r[53];
assign temp_mult[822] = 16'd1390 * d1_input_r[54];
assign temp_mult[823] = 16'd1097 * d1_input_r[55];
assign temp_mult[824] = 16'd1419 * d1_input_r[56];
assign temp_mult[825] = 16'd35001 * d1_input_r[57];
assign temp_mult[826] = 16'd3022 * d1_input_r[58];
assign temp_mult[827] = 16'd35292 * d1_input_r[59];
assign temp_mult[828] = 16'd35208 * d1_input_r[60];
assign temp_mult[829] = 16'd34584 * d1_input_r[61];
assign temp_mult[830] = 16'd2189 * d1_input_r[62];
assign temp_mult[831] = 16'd33479 * d1_input_r[63];
assign temp_mult[832] = 16'd35315 * d1_input_r[64];
assign temp_mult[833] = 16'd836 * d1_input_r[65];
assign temp_mult[834] = 16'd2041 * d1_input_r[66];
assign temp_mult[835] = 16'd35457 * d1_input_r[67];
assign temp_mult[836] = 16'd1651 * d1_input_r[68];
assign temp_mult[837] = 16'd828 * d1_input_r[69];
assign temp_mult[838] = 16'd872 * d1_input_r[70];
assign temp_mult[839] = 16'd539 * d1_input_r[71];
assign temp_mult[840] = 16'd1319 * d1_input_r[72];
assign temp_mult[841] = 16'd34557 * d1_input_r[73];
assign temp_mult[842] = 16'd33301 * d1_input_r[74];
assign temp_mult[843] = 16'd579 * d1_input_r[75];
assign temp_mult[844] = 16'd33173 * d1_input_r[76];
assign temp_mult[845] = 16'd334 * d1_input_r[77];
assign temp_mult[846] = 16'd2210 * d1_input_r[78];
assign temp_mult[847] = 16'd2884 * d1_input_r[79];
assign temp_mult[848] = 16'd1616 * d1_input_r[80];
assign temp_mult[849] = 16'd33196 * d1_input_r[81];
assign temp_mult[850] = 16'd873 * d1_input_r[82];
assign temp_mult[851] = 16'd33970 * d1_input_r[83];
assign temp_mult[852] = 16'd1410 * d1_input_r[84];
assign temp_mult[853] = 16'd34550 * d1_input_r[85];
assign temp_mult[854] = 16'd34430 * d1_input_r[86];
assign temp_mult[855] = 16'd33926 * d1_input_r[87];
assign temp_mult[856] = 16'd35229 * d1_input_r[88];
assign temp_mult[857] = 16'd2849 * d1_input_r[89];
assign temp_mult[858] = 16'd801 * d1_input_r[90];
assign temp_mult[859] = 16'd34141 * d1_input_r[91];
assign temp_mult[860] = 16'd33958 * d1_input_r[92];
assign temp_mult[861] = 16'd2924 * d1_input_r[93];
assign temp_mult[862] = 16'd1920 * d1_input_r[94];
assign temp_mult[863] = 16'd35771 * d1_input_r[95];
assign temp_mult[864] = 16'd1843 * d1_input_r[96];
assign temp_mult[865] = 16'd513 * d1_input_r[97];
assign temp_mult[866] = 16'd33657 * d1_input_r[98];
assign temp_mult[867] = 16'd35732 * d1_input_r[99];
assign temp_mult[868] = 16'd2142 * d1_input_r[100];
assign temp_mult[869] = 16'd2260 * d1_input_r[101];
assign temp_mult[870] = 16'd2037 * d1_input_r[102];
assign temp_mult[871] = 16'd33969 * d1_input_r[103];
assign temp_mult[872] = 16'd35041 * d1_input_r[104];
assign temp_mult[873] = 16'd2275 * d1_input_r[105];
assign temp_mult[874] = 16'd354 * d1_input_r[106];
assign temp_mult[875] = 16'd34734 * d1_input_r[107];
assign temp_mult[876] = 16'd122 * d1_input_r[108];
assign temp_mult[877] = 16'd1517 * d1_input_r[109];
assign temp_mult[878] = 16'd1969 * d1_input_r[110];
assign temp_mult[879] = 16'd32775 * d1_input_r[111];
assign temp_mult[880] = 16'd33170 * d1_input_r[112];
assign temp_mult[881] = 16'd34598 * d1_input_r[113];
assign temp_mult[882] = 16'd34679 * d1_input_r[114];
assign temp_mult[883] = 16'd33162 * d1_input_r[115];
assign temp_mult[884] = 16'd554 * d1_input_r[116];
assign temp_mult[885] = 16'd34034 * d1_input_r[117];
assign temp_mult[886] = 16'd33987 * d1_input_r[118];
assign temp_mult[887] = 16'd1250 * d1_input_r[119];
assign temp_mult[888] = 16'd32908 * d1_input_r[120];
assign temp_mult[889] = 16'd33551 * d1_input_r[121];
assign temp_mult[890] = 16'd1151 * d1_input_r[122];
assign temp_mult[891] = 16'd35741 * d1_input_r[123];
assign temp_mult[892] = 16'd1221 * d1_input_r[124];
assign temp_mult[893] = 16'd34138 * d1_input_r[125];
assign temp_mult[894] = 16'd1526 * d1_input_r[126];
assign temp_mult[895] = 16'd1135 * d1_input_r[127];
assign temp_mult[896] = 16'd35909 * d1_input_r[128];
assign temp_mult[897] = 16'd1661 * d1_input_r[129];
assign temp_mult[898] = 16'd33812 * d1_input_r[130];
assign temp_mult[899] = 16'd34957 * d1_input_r[131];
assign temp_mult[900] = 16'd2074 * d1_input_r[132];
assign temp_mult[901] = 16'd1265 * d1_input_r[133];
assign temp_mult[902] = 16'd1475 * d1_input_r[134];
assign temp_mult[903] = 16'd1647 * d1_input_r[135];
assign temp_mult[904] = 16'd447 * d1_input_r[136];
assign temp_mult[905] = 16'd33853 * d1_input_r[137];
assign temp_mult[906] = 16'd2479 * d1_input_r[138];
assign temp_mult[907] = 16'd486 * d1_input_r[139];
assign temp_mult[908] = 16'd33967 * d1_input_r[140];
assign temp_mult[909] = 16'd33295 * d1_input_r[141];
assign temp_mult[910] = 16'd34128 * d1_input_r[142];
assign temp_mult[911] = 16'd994 * d1_input_r[143];
assign temp_mult[912] = 16'd2530 * d1_input_r[144];
assign temp_mult[913] = 16'd33961 * d1_input_r[145];
assign temp_mult[914] = 16'd34945 * d1_input_r[146];
assign temp_mult[915] = 16'd34327 * d1_input_r[147];
assign temp_mult[916] = 16'd2964 * d1_input_r[148];
assign temp_mult[917] = 16'd1666 * d1_input_r[149];
assign temp_mult[918] = 16'd1429 * d1_input_r[150];
assign temp_mult[919] = 16'd33167 * d1_input_r[151];
assign temp_mult[920] = 16'd34985 * d1_input_r[152];
assign temp_mult[921] = 16'd2347 * d1_input_r[153];
assign temp_mult[922] = 16'd33469 * d1_input_r[154];
assign temp_mult[923] = 16'd32852 * d1_input_r[155];
assign temp_mult[924] = 16'd222 * d1_input_r[156];
assign temp_mult[925] = 16'd2049 * d1_input_r[157];
assign temp_mult[926] = 16'd1790 * d1_input_r[158];
assign temp_mult[927] = 16'd680 * d1_input_r[159];
assign temp_mult[928] = 16'd34420 * d1_input_r[160];
assign temp_mult[929] = 16'd2229 * d1_input_r[161];
assign temp_mult[930] = 16'd679 * d1_input_r[162];
assign temp_mult[931] = 16'd1516 * d1_input_r[163];
assign temp_mult[932] = 16'd1727 * d1_input_r[164];
assign temp_mult[933] = 16'd2135 * d1_input_r[165];
assign temp_mult[934] = 16'd34397 * d1_input_r[166];
assign temp_mult[935] = 16'd33511 * d1_input_r[167];
assign temp_mult[936] = 16'd1000 * d1_input_r[168];
assign temp_mult[937] = 16'd33422 * d1_input_r[169];
assign temp_mult[938] = 16'd705 * d1_input_r[170];
assign temp_mult[939] = 16'd1811 * d1_input_r[171];
assign temp_mult[940] = 16'd33699 * d1_input_r[172];
assign temp_mult[941] = 16'd397 * d1_input_r[173];
assign temp_mult[942] = 16'd33596 * d1_input_r[174];
assign temp_mult[943] = 16'd433 * d1_input_r[175];
assign temp_mult[944] = 16'd33237 * d1_input_r[176];
assign temp_mult[945] = 16'd33933 * d1_input_r[177];
assign temp_mult[946] = 16'd34933 * d1_input_r[178];
assign temp_mult[947] = 16'd34687 * d1_input_r[179];
assign temp_mult[948] = 16'd2713 * d1_input_r[180];
assign temp_mult[949] = 16'd1122 * d1_input_r[181];
assign temp_mult[950] = 16'd33737 * d1_input_r[182];
assign temp_mult[951] = 16'd33743 * d1_input_r[183];
assign temp_mult[952] = 16'd793 * d1_input_r[184];
assign temp_mult[953] = 16'd2496 * d1_input_r[185];
assign temp_mult[954] = 16'd33328 * d1_input_r[186];
assign temp_mult[955] = 16'd803 * d1_input_r[187];
assign temp_mult[956] = 16'd33001 * d1_input_r[188];
assign temp_mult[957] = 16'd2735 * d1_input_r[189];
assign temp_mult[958] = 16'd1950 * d1_input_r[190];
assign temp_mult[959] = 16'd535 * d1_input_r[191];
assign temp_mult[960] = 16'd35031 * d1_input_r[192];
assign temp_mult[961] = 16'd1216 * d1_input_r[193];
assign temp_mult[962] = 16'd34730 * d1_input_r[194];
assign temp_mult[963] = 16'd32871 * d1_input_r[195];
assign temp_mult[964] = 16'd802 * d1_input_r[196];
assign temp_mult[965] = 16'd662 * d1_input_r[197];
assign temp_mult[966] = 16'd33743 * d1_input_r[198];
assign temp_mult[967] = 16'd516 * d1_input_r[199];
assign temp_mult[968] = 16'd35665 * d1_input_r[200];
assign temp_mult[969] = 16'd774 * d1_input_r[201];
assign temp_mult[970] = 16'd939 * d1_input_r[202];
assign temp_mult[971] = 16'd32816 * d1_input_r[203];
assign temp_mult[972] = 16'd34150 * d1_input_r[204];
assign temp_mult[973] = 16'd35420 * d1_input_r[205];
assign temp_mult[974] = 16'd1456 * d1_input_r[206];
assign temp_mult[975] = 16'd501 * d1_input_r[207];
assign temp_mult[976] = 16'd1190 * d1_input_r[208];
assign temp_mult[977] = 16'd34887 * d1_input_r[209];
assign temp_mult[978] = 16'd32966 * d1_input_r[210];
assign temp_mult[979] = 16'd34150 * d1_input_r[211];
assign temp_mult[980] = 16'd3008 * d1_input_r[212];
assign temp_mult[981] = 16'd34244 * d1_input_r[213];
assign temp_mult[982] = 16'd33623 * d1_input_r[214];
assign temp_mult[983] = 16'd1685 * d1_input_r[215];
assign temp_mult[984] = 16'd33213 * d1_input_r[216];
assign temp_mult[985] = 16'd2179 * d1_input_r[217];
assign temp_mult[986] = 16'd34125 * d1_input_r[218];
assign temp_mult[987] = 16'd1115 * d1_input_r[219];
assign temp_mult[988] = 16'd33935 * d1_input_r[220];
assign temp_mult[989] = 16'd2460 * d1_input_r[221];
assign temp_mult[990] = 16'd33038 * d1_input_r[222];
assign temp_mult[991] = 16'd33541 * d1_input_r[223];
assign temp_mult[992] = 16'd33742 * d1_input_r[224];
assign temp_mult[993] = 16'd1472 * d1_input_r[225];
assign temp_mult[994] = 16'd33436 * d1_input_r[226];
assign temp_mult[995] = 16'd1044 * d1_input_r[227];
assign temp_mult[996] = 16'd705 * d1_input_r[228];
assign temp_mult[997] = 16'd33431 * d1_input_r[229];
assign temp_mult[998] = 16'd34594 * d1_input_r[230];
assign temp_mult[999] = 16'd33268 * d1_input_r[231];
assign temp_mult[1000] = 16'd34076 * d1_input_r[232];
assign temp_mult[1001] = 16'd1060 * d1_input_r[233];
assign temp_mult[1002] = 16'd32906 * d1_input_r[234];
assign temp_mult[1003] = 16'd34681 * d1_input_r[235];
assign temp_mult[1004] = 16'd33523 * d1_input_r[236];
assign temp_mult[1005] = 16'd34134 * d1_input_r[237];
assign temp_mult[1006] = 16'd1900 * d1_input_r[238];
assign temp_mult[1007] = 16'd2208 * d1_input_r[239];
assign temp_mult[1008] = 16'd1292 * d1_input_r[240];
assign temp_mult[1009] = 16'd1152 * d1_input_r[241];
assign temp_mult[1010] = 16'd35077 * d1_input_r[242];
assign temp_mult[1011] = 16'd33308 * d1_input_r[243];
assign temp_mult[1012] = 16'd34095 * d1_input_r[244];
assign temp_mult[1013] = 16'd2222 * d1_input_r[245];
assign temp_mult[1014] = 16'd34935 * d1_input_r[246];
assign temp_mult[1015] = 16'd34745 * d1_input_r[247];
assign temp_mult[1016] = 16'd34674 * d1_input_r[248];
assign temp_mult[1017] = 16'd2328 * d1_input_r[249];
assign temp_mult[1018] = 16'd34186 * d1_input_r[250];
assign temp_mult[1019] = 16'd34893 * d1_input_r[251];
assign temp_mult[1020] = 16'd35358 * d1_input_r[252];
assign temp_mult[1021] = 16'd33389 * d1_input_r[253];
assign temp_mult[1022] = 16'd291 * d1_input_r[254];
assign temp_mult[1023] = 16'd35035 * d1_input_r[255];


always @(*) begin
	if(!rst_n) begin
		for(j = 0; j < 256; j = j+1) begin
			d1_input_r[j] = 16'd0;
		end
	end
	else begin
		for(j = 0; j < 256; j = j+1) begin
			d1_input_r[j] = d1_input[((16*(j+1))-1) -: 16];
		end
	end
end


always @(*) begin
	if(!rst_n) begin
		temp_add[0] = 16'd0;
		temp_add[1] = 16'd0;
		temp_add[2] = 16'd0;
		temp_add[3] = 16'd0;
	end
	else begin
		for(i = 0; i < 256; i = i+1) begin
			temp_add[0] = temp_add[0] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
		for(i = 256; i < 512; i = i+1) begin
			temp_add[1] = temp_add[1] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
		for(i = 512; i < 768; i = i+1) begin
			temp_add[2] = temp_add[2] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
		for(i = 768; i < 1024; i = i+1) begin
			temp_add[3] = temp_add[3] + {temp_mult[i][31], temp_mult[i][29], temp_mult[i][27:14]};
		end
	end
end

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		d1_output <= 64'd0;
	end
	else begin
		d1_output[15:0] <= temp_add[0] + bias[0];
		d1_output[31:16] <= temp_add[1] + bias[1];
		d1_output[47:32] <= temp_add[2] + bias[2];
		d1_output[63:48] <= temp_add[3] + bias[3];
	end
end

endmodule